/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Nov  5 21:59:42 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1099544531 */

module addition_normaliser(in_e, in_m, out_e, out_m);
   input [7:0]in_e;
   input [24:0]in_m;
   output [7:0]out_e;
   output [24:0]out_m;

   wire n_0_23;
   wire n_0_2;
   wire n_0_24;
   wire n_0_1;
   wire n_0_25;
   wire n_0_0;
   wire n_0_26;
   wire n_0_3;
   wire n_0_27;
   wire n_0_4;
   wire n_0_28;
   wire n_0_5;
   wire n_0_29;
   wire n_0_6;
   wire n_0_30;
   wire n_0_7;
   wire n_0_31;
   wire n_0_8;
   wire n_0_32;
   wire n_0_9;
   wire n_0_33;
   wire n_0_10;
   wire n_0_34;
   wire n_0_11;
   wire n_0_35;
   wire n_0_12;
   wire n_0_36;
   wire n_0_13;
   wire n_0_37;
   wire n_0_14;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_15;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_16;
   wire n_0_17;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_18;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_19;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_20;
   wire n_0_186;
   wire n_0_21;
   wire n_0_187;
   wire n_0_188;
   wire n_0_22;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_317;
   wire n_0_318;
   wire n_0_319;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_332;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_337;
   wire n_0_338;
   wire n_0_339;
   wire n_0_340;
   wire n_0_341;
   wire n_0_342;
   wire n_0_343;
   wire n_0_344;
   wire n_0_345;
   wire n_0_346;
   wire n_0_347;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_355;
   wire n_0_356;
   wire n_0_357;
   wire n_0_358;
   wire n_0_359;
   wire n_0_360;
   wire n_0_361;
   wire n_0_362;
   wire n_0_363;
   wire n_0_364;
   wire n_0_365;
   wire n_0_366;
   wire n_0_367;
   wire n_0_368;
   wire n_0_369;
   wire n_0_370;
   wire n_0_371;
   wire n_0_372;
   wire n_0_373;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_377;
   wire n_0_378;
   wire n_0_379;
   wire n_0_380;
   wire n_0_381;
   wire n_0_382;
   wire n_0_383;
   wire n_0_384;
   wire n_0_385;
   wire n_0_386;
   wire n_0_387;
   wire n_0_388;
   wire n_0_389;
   wire n_0_390;
   wire n_0_391;
   wire n_0_392;
   wire n_0_393;
   wire n_0_394;
   wire n_0_395;
   wire n_0_396;
   wire n_0_397;
   wire n_0_398;
   wire n_0_399;
   wire n_0_400;
   wire n_0_401;
   wire n_0_402;
   wire n_0_403;
   wire n_0_404;
   wire n_0_405;
   wire n_0_406;
   wire n_0_407;
   wire n_0_408;
   wire n_0_409;
   wire n_0_410;
   wire n_0_411;
   wire n_0_412;
   wire n_0_413;
   wire n_0_414;
   wire n_0_415;
   wire n_0_416;
   wire n_0_417;
   wire n_0_418;
   wire n_0_419;
   wire n_0_420;
   wire n_0_421;
   wire n_0_422;
   wire n_0_423;
   wire n_0_424;
   wire n_0_425;
   wire n_0_426;
   wire n_0_427;
   wire n_0_428;
   wire n_0_429;
   wire n_0_430;
   wire n_0_431;
   wire n_0_432;
   wire n_0_433;
   wire n_0_434;
   wire n_0_435;
   wire n_0_436;
   wire n_0_437;
   wire n_0_438;
   wire n_0_439;
   wire n_0_440;
   wire n_0_441;
   wire n_0_442;
   wire n_0_443;
   wire n_0_444;
   wire n_0_445;
   wire n_0_446;
   wire n_0_447;
   wire n_0_448;
   wire n_0_449;
   wire n_0_450;
   wire n_0_451;
   wire n_0_452;
   wire n_0_453;
   wire n_0_454;
   wire n_0_455;
   wire n_0_456;
   wire n_0_457;
   wire n_0_458;
   wire n_0_459;
   wire n_0_460;
   wire n_0_461;
   wire n_0_462;
   wire n_0_463;
   wire n_0_464;
   wire n_0_465;
   wire n_0_466;
   wire n_0_467;
   wire n_0_468;
   wire n_0_469;
   wire n_0_470;
   wire n_0_471;
   wire n_0_472;
   wire n_0_473;
   wire n_0_474;
   wire n_0_475;
   wire n_0_476;
   wire n_0_477;
   wire n_0_478;
   wire n_0_479;
   wire n_0_480;
   wire n_0_481;
   wire n_0_482;
   wire n_0_483;
   wire n_0_484;
   wire n_0_485;
   wire n_0_486;
   wire n_0_487;
   wire n_0_488;
   wire n_0_489;
   wire n_0_490;
   wire n_0_491;
   wire n_0_492;
   wire n_0_493;
   wire n_0_494;
   wire n_0_495;
   wire n_0_496;
   wire n_0_497;
   wire n_0_498;
   wire n_0_499;
   wire n_0_500;
   wire n_0_501;
   wire n_0_502;
   wire n_0_503;
   wire n_0_504;
   wire n_0_505;
   wire n_0_506;
   wire n_0_507;
   wire n_0_508;
   wire n_0_509;
   wire n_0_510;
   wire n_0_511;
   wire n_0_512;
   wire n_0_513;
   wire n_0_514;

   DLH_X1 \out_m_reg[22]  (.D(n_30), .G(n_8), .Q(out_m[22]));
   DLH_X1 \out_m_reg[21]  (.D(n_29), .G(n_8), .Q(out_m[21]));
   DLH_X1 \out_m_reg[20]  (.D(n_28), .G(n_8), .Q(out_m[20]));
   DLH_X1 \out_m_reg[19]  (.D(n_27), .G(n_8), .Q(out_m[19]));
   DLH_X1 \out_m_reg[18]  (.D(n_26), .G(n_8), .Q(out_m[18]));
   DLH_X1 \out_m_reg[17]  (.D(n_25), .G(n_8), .Q(out_m[17]));
   DLH_X1 \out_m_reg[16]  (.D(n_24), .G(n_8), .Q(out_m[16]));
   DLH_X1 \out_m_reg[15]  (.D(n_23), .G(n_8), .Q(out_m[15]));
   DLH_X1 \out_m_reg[14]  (.D(n_22), .G(n_8), .Q(out_m[14]));
   DLH_X1 \out_m_reg[13]  (.D(n_21), .G(n_8), .Q(out_m[13]));
   DLH_X1 \out_m_reg[12]  (.D(n_20), .G(n_8), .Q(out_m[12]));
   DLH_X1 \out_m_reg[11]  (.D(n_19), .G(n_8), .Q(out_m[11]));
   DLH_X1 \out_m_reg[10]  (.D(n_18), .G(n_8), .Q(out_m[10]));
   DLH_X1 \out_m_reg[9]  (.D(n_17), .G(n_8), .Q(out_m[9]));
   DLH_X1 \out_m_reg[8]  (.D(n_16), .G(n_8), .Q(out_m[8]));
   DLH_X1 \out_m_reg[7]  (.D(n_15), .G(n_8), .Q(out_m[7]));
   DLH_X1 \out_m_reg[6]  (.D(n_14), .G(n_8), .Q(out_m[6]));
   DLH_X1 \out_m_reg[5]  (.D(n_13), .G(n_8), .Q(out_m[5]));
   DLH_X1 \out_m_reg[4]  (.D(n_12), .G(n_8), .Q(out_m[4]));
   DLH_X1 \out_m_reg[3]  (.D(n_11), .G(n_8), .Q(out_m[3]));
   DLH_X1 \out_m_reg[2]  (.D(n_10), .G(n_8), .Q(out_m[2]));
   DLH_X1 \out_m_reg[1]  (.D(n_9), .G(n_8), .Q(out_m[1]));
   DLH_X1 \out_e_reg[7]  (.D(n_7), .G(n_8), .Q(out_e[7]));
   DLH_X1 \out_e_reg[6]  (.D(n_6), .G(n_8), .Q(out_e[6]));
   DLH_X1 \out_e_reg[5]  (.D(n_5), .G(n_8), .Q(out_e[5]));
   DLH_X1 \out_e_reg[4]  (.D(n_4), .G(n_8), .Q(out_e[4]));
   DLH_X1 \out_e_reg[3]  (.D(n_3), .G(n_8), .Q(out_e[3]));
   DLH_X1 \out_e_reg[2]  (.D(n_2), .G(n_8), .Q(out_e[2]));
   DLH_X1 \out_e_reg[1]  (.D(n_1), .G(n_8), .Q(out_e[1]));
   DLH_X1 \out_e_reg[0]  (.D(n_0), .G(n_8), .Q(out_e[0]));
   HA_X1 i_0_0 (.A(in_e[3]), .B(n_0_20), .CO(n_0_2), .S(n_0_23));
   HA_X1 i_0_1 (.A(in_e[3]), .B(n_0_22), .CO(n_0_1), .S(n_0_24));
   HA_X1 i_0_2 (.A(in_e[3]), .B(n_0_19), .CO(n_0_0), .S(n_0_25));
   HA_X1 i_0_3 (.A(in_e[3]), .B(in_e[2]), .CO(n_0_3), .S(n_0_26));
   HA_X1 i_0_4 (.A(in_e[3]), .B(n_0_12), .CO(n_0_4), .S(n_0_27));
   HA_X1 i_0_5 (.A(in_e[3]), .B(n_0_13), .CO(n_0_5), .S(n_0_28));
   HA_X1 i_0_6 (.A(in_e[3]), .B(n_0_14), .CO(n_0_6), .S(n_0_29));
   HA_X1 i_0_7 (.A(in_e[4]), .B(n_0_16), .CO(n_0_7), .S(n_0_30));
   HA_X1 i_0_8 (.A(in_e[4]), .B(n_0_17), .CO(n_0_8), .S(n_0_31));
   HA_X1 i_0_9 (.A(in_e[4]), .B(n_0_15), .CO(n_0_9), .S(n_0_32));
   HA_X1 i_0_10 (.A(in_e[4]), .B(n_0_18), .CO(n_0_10), .S(n_0_33));
   HA_X1 i_0_11 (.A(in_e[1]), .B(in_e[0]), .CO(n_0_11), .S(n_0_34));
   HA_X1 i_0_12 (.A(in_e[2]), .B(n_0_21), .CO(n_0_12), .S(n_0_35));
   HA_X1 i_0_13 (.A(in_e[2]), .B(in_e[1]), .CO(n_0_13), .S(n_0_36));
   HA_X1 i_0_14 (.A(in_e[2]), .B(n_0_11), .CO(n_0_14), .S(n_0_37));
   XOR2_X1 i_0_15 (.A(in_e[0]), .B(n_0_38), .Z(n_0));
   AOI221_X1 i_0_16 (.A(n_0_353), .B1(n_0_403), .B2(n_0_402), .C1(n_0_166), 
      .C2(n_0_39), .ZN(n_0_38));
   OAI211_X1 i_0_17 (.A(n_0_503), .B(n_0_361), .C1(n_0_467), .C2(n_0_40), 
      .ZN(n_0_39));
   AOI21_X1 i_0_18 (.A(in_m[11]), .B1(n_0_334), .B2(n_0_41), .ZN(n_0_40));
   AOI21_X1 i_0_19 (.A(in_m[10]), .B1(n_0_161), .B2(n_0_42), .ZN(n_0_41));
   NOR3_X1 i_0_20 (.A1(in_m[9]), .A2(in_m[7]), .A3(n_0_433), .ZN(n_0_42));
   NAND4_X1 i_0_21 (.A1(n_0_68), .A2(n_0_53), .A3(n_0_43), .A4(n_0_47), .ZN(n_1));
   INV_X1 i_0_22 (.A(n_0_44), .ZN(n_0_43));
   AOI211_X1 i_0_23 (.A(n_0_165), .B(n_0_74), .C1(n_0_501), .C2(n_0_45), 
      .ZN(n_0_44));
   NAND2_X1 i_0_24 (.A1(n_0_453), .A2(n_0_46), .ZN(n_0_45));
   AOI22_X1 i_0_25 (.A1(n_0_51), .A2(n_0_48), .B1(in_m[10]), .B2(n_0_76), 
      .ZN(n_0_46));
   AOI221_X1 i_0_26 (.A(n_0_60), .B1(in_e[1]), .B2(n_0_77), .C1(n_0_34), 
      .C2(n_0_64), .ZN(n_0_47));
   AOI21_X1 i_0_27 (.A(n_0_448), .B1(n_0_34), .B2(n_0_49), .ZN(n_0_48));
   NAND2_X1 i_0_28 (.A1(n_0_496), .A2(n_0_50), .ZN(n_0_49));
   NAND3_X1 i_0_29 (.A1(n_0_495), .A2(in_m[4]), .A3(n_0_494), .ZN(n_0_50));
   NAND2_X1 i_0_30 (.A1(n_0_496), .A2(n_0_52), .ZN(n_0_51));
   AOI21_X1 i_0_31 (.A(in_m[7]), .B1(n_0_434), .B2(n_0_59), .ZN(n_0_52));
   NAND3_X1 i_0_32 (.A1(n_0_166), .A2(n_0_70), .A3(n_0_54), .ZN(n_0_53));
   OAI221_X1 i_0_33 (.A(n_0_503), .B1(n_0_76), .B2(n_0_63), .C1(n_0_425), 
      .C2(n_0_55), .ZN(n_0_54));
   AOI221_X1 i_0_34 (.A(n_0_56), .B1(n_0_34), .B2(n_0_57), .C1(n_0_329), 
      .C2(n_0_58), .ZN(n_0_55));
   OAI21_X1 i_0_35 (.A(n_0_499), .B1(n_0_498), .B2(n_0_76), .ZN(n_0_56));
   AOI21_X1 i_0_36 (.A(n_0_448), .B1(n_0_496), .B2(n_0_157), .ZN(n_0_57));
   NAND3_X1 i_0_37 (.A1(n_0_495), .A2(n_0_161), .A3(n_0_59), .ZN(n_0_58));
   NAND2_X1 i_0_38 (.A1(in_m[6]), .A2(n_0_75), .ZN(n_0_59));
   AOI211_X1 i_0_39 (.A(in_e[1]), .B(n_0_483), .C1(n_0_509), .C2(n_0_61), 
      .ZN(n_0_60));
   NAND3_X1 i_0_40 (.A1(n_0_508), .A2(n_0_507), .A3(n_0_62), .ZN(n_0_61));
   OAI22_X1 i_0_41 (.A1(in_m[18]), .A2(n_0_505), .B1(n_0_76), .B2(n_0_63), 
      .ZN(n_0_62));
   AOI21_X1 i_0_42 (.A(in_m[18]), .B1(in_m[14]), .B2(n_0_469), .ZN(n_0_63));
   OR2_X1 i_0_43 (.A1(n_0_351), .A2(n_0_65), .ZN(n_0_64));
   OAI33_X1 i_0_44 (.A1(n_0_500), .A2(n_0_165), .A3(n_0_67), .B1(n_0_504), 
      .B2(n_0_324), .B3(n_0_66), .ZN(n_0_65));
   AOI21_X1 i_0_45 (.A(n_0_70), .B1(n_0_511), .B2(n_0_507), .ZN(n_0_66));
   AOI21_X1 i_0_46 (.A(n_0_73), .B1(n_0_501), .B2(n_0_70), .ZN(n_0_67));
   OAI21_X1 i_0_47 (.A(n_0_75), .B1(n_0_483), .B2(n_0_69), .ZN(n_0_68));
   OAI33_X1 i_0_48 (.A1(n_0_363), .A2(n_0_72), .A3(n_0_191), .B1(in_m[13]), 
      .B2(n_0_71), .B3(n_0_199), .ZN(n_0_69));
   INV_X1 i_0_49 (.A(n_0_71), .ZN(n_0_70));
   NAND3_X1 i_0_50 (.A1(in_e[1]), .A2(n_0_509), .A3(n_0_505), .ZN(n_0_71));
   NAND3_X1 i_0_51 (.A1(n_0_496), .A2(n_0_458), .A3(n_0_73), .ZN(n_0_72));
   INV_X1 i_0_52 (.A(n_0_74), .ZN(n_0_73));
   NAND3_X1 i_0_53 (.A1(n_0_511), .A2(n_0_507), .A3(n_0_503), .ZN(n_0_74));
   INV_X1 i_0_54 (.A(n_0_76), .ZN(n_0_75));
   AOI21_X1 i_0_55 (.A(n_0_186), .B1(in_e[1]), .B2(in_e[0]), .ZN(n_0_76));
   OAI22_X1 i_0_56 (.A1(n_0_507), .A2(n_0_478), .B1(n_0_510), .B2(n_0_308), 
      .ZN(n_0_77));
   NAND4_X1 i_0_57 (.A1(n_0_89), .A2(n_0_81), .A3(n_0_78), .A4(n_0_90), .ZN(n_2));
   AOI22_X1 i_0_58 (.A1(n_0_164), .A2(n_0_80), .B1(n_0_103), .B2(n_0_79), 
      .ZN(n_0_78));
   AOI211_X1 i_0_59 (.A(n_0_165), .B(n_0_453), .C1(in_m[12]), .C2(n_0_97), 
      .ZN(n_0_79));
   AOI22_X1 i_0_60 (.A1(n_0_83), .A2(n_0_82), .B1(n_0_106), .B2(n_0_104), 
      .ZN(n_0_80));
   AOI222_X1 i_0_61 (.A1(n_0_37), .A2(n_0_322), .B1(n_0_36), .B2(n_0_310), 
      .C1(n_0_351), .C2(n_0_96), .ZN(n_0_81));
   AOI21_X1 i_0_62 (.A(n_0_84), .B1(n_0_37), .B2(n_0_333), .ZN(n_0_82));
   AOI22_X1 i_0_63 (.A1(in_m[10]), .A2(n_0_35), .B1(n_0_36), .B2(n_0_422), 
      .ZN(n_0_83));
   AOI221_X1 i_0_64 (.A(n_0_330), .B1(in_m[7]), .B2(n_0_106), .C1(n_0_86), 
      .C2(n_0_85), .ZN(n_0_84));
   AOI221_X1 i_0_65 (.A(in_m[7]), .B1(n_0_156), .B2(n_0_96), .C1(n_0_160), 
      .C2(n_0_103), .ZN(n_0_85));
   OAI211_X1 i_0_66 (.A(n_0_87), .B(n_0_394), .C1(in_e[2]), .C2(n_0_88), 
      .ZN(n_0_86));
   NAND2_X1 i_0_67 (.A1(in_e[2]), .A2(n_0_88), .ZN(n_0_87));
   OAI21_X1 i_0_68 (.A(n_0_21), .B1(in_e[1]), .B2(in_m[6]), .ZN(n_0_88));
   AOI22_X1 i_0_69 (.A1(n_0_404), .A2(n_0_188), .B1(n_0_35), .B2(n_0_309), 
      .ZN(n_0_89));
   AOI22_X1 i_0_70 (.A1(n_0_108), .A2(n_0_100), .B1(n_0_92), .B2(n_0_91), 
      .ZN(n_0_90));
   NAND2_X1 i_0_71 (.A1(in_e[2]), .A2(n_0_93), .ZN(n_0_91));
   OAI221_X1 i_0_72 (.A(n_0_512), .B1(n_0_507), .B2(n_0_478), .C1(n_0_290), 
      .C2(n_0_98), .ZN(n_0_92));
   AOI22_X1 i_0_73 (.A1(in_e[1]), .A2(n_0_404), .B1(n_0_415), .B2(n_0_94), 
      .ZN(n_0_93));
   OAI21_X1 i_0_74 (.A(n_0_503), .B1(n_0_99), .B2(n_0_95), .ZN(n_0_94));
   AOI21_X1 i_0_75 (.A(n_0_455), .B1(in_m[12]), .B2(n_0_96), .ZN(n_0_95));
   INV_X1 i_0_76 (.A(n_0_97), .ZN(n_0_96));
   AOI21_X1 i_0_77 (.A(n_0_181), .B1(in_e[2]), .B2(n_0_11), .ZN(n_0_97));
   INV_X1 i_0_78 (.A(n_0_99), .ZN(n_0_98));
   AOI211_X1 i_0_79 (.A(in_e[1]), .B(n_0_454), .C1(in_e[0]), .C2(in_m[14]), 
      .ZN(n_0_99));
   OAI21_X1 i_0_80 (.A(n_0_101), .B1(n_0_199), .B2(n_0_102), .ZN(n_0_100));
   AOI21_X1 i_0_81 (.A(n_0_483), .B1(n_0_198), .B2(n_0_107), .ZN(n_0_101));
   NAND2_X1 i_0_82 (.A1(n_0_495), .A2(n_0_103), .ZN(n_0_102));
   INV_X1 i_0_83 (.A(n_0_104), .ZN(n_0_103));
   NAND3_X1 i_0_84 (.A1(n_0_512), .A2(n_0_509), .A3(n_0_105), .ZN(n_0_104));
   NOR3_X1 i_0_85 (.A1(in_m[17]), .A2(in_m[15]), .A3(in_m[13]), .ZN(n_0_105));
   INV_X1 i_0_86 (.A(n_0_107), .ZN(n_0_106));
   NOR2_X1 i_0_87 (.A1(n_0_512), .A2(n_0_197), .ZN(n_0_107));
   OAI21_X1 i_0_88 (.A(n_0_20), .B1(n_0_512), .B2(n_0_186), .ZN(n_0_108));
   OAI221_X1 i_0_89 (.A(n_0_109), .B1(n_0_128), .B2(n_0_126), .C1(in_e[3]), 
      .C2(n_0_179), .ZN(n_3));
   AOI21_X1 i_0_90 (.A(n_0_110), .B1(in_e[3]), .B2(n_0_129), .ZN(n_0_109));
   INV_X1 i_0_91 (.A(n_0_111), .ZN(n_0_110));
   AOI211_X1 i_0_92 (.A(n_0_115), .B(n_0_114), .C1(n_0_163), .C2(n_0_112), 
      .ZN(n_0_111));
   AOI211_X1 i_0_93 (.A(n_0_124), .B(n_0_113), .C1(in_m[6]), .C2(n_0_128), 
      .ZN(n_0_112));
   OAI221_X1 i_0_94 (.A(n_0_127), .B1(n_0_434), .B2(n_0_125), .C1(n_0_394), 
      .C2(n_0_122), .ZN(n_0_113));
   OAI211_X1 i_0_95 (.A(n_0_116), .B(n_0_118), .C1(n_0_352), .C2(n_0_15), 
      .ZN(n_0_114));
   OAI33_X1 i_0_96 (.A1(n_0_334), .A2(n_0_175), .A3(n_0_486), .B1(n_0_416), 
      .B2(n_0_297), .B3(n_0_117), .ZN(n_0_115));
   NAND2_X1 i_0_97 (.A1(n_0_513), .A2(n_0_181), .ZN(n_0_15));
   NAND2_X1 i_0_98 (.A1(n_0_404), .A2(n_0_125), .ZN(n_0_116));
   NAND2_X1 i_0_99 (.A1(n_0_503), .A2(n_0_28), .ZN(n_0_117));
   INV_X1 i_0_100 (.A(n_0_119), .ZN(n_0_118));
   AOI21_X1 i_0_101 (.A(n_0_436), .B1(n_0_121), .B2(n_0_120), .ZN(n_0_119));
   AOI22_X1 i_0_102 (.A1(n_0_26), .A2(n_0_347), .B1(n_0_27), .B2(n_0_315), 
      .ZN(n_0_120));
   AOI222_X1 i_0_103 (.A1(in_m[14]), .A2(n_0_23), .B1(n_0_24), .B2(n_0_360), 
      .C1(n_0_25), .C2(n_0_383), .ZN(n_0_121));
   AOI22_X1 i_0_104 (.A1(n_0_492), .A2(n_0_491), .B1(n_0_18), .B2(n_0_123), 
      .ZN(n_0_122));
   OAI211_X1 i_0_105 (.A(in_e[3]), .B(n_0_19), .C1(in_e[2]), .C2(in_m[4]), 
      .ZN(n_0_123));
   AND3_X1 i_0_106 (.A1(n_0_513), .A2(n_0_11), .A3(n_0_156), .ZN(n_0_124));
   OAI21_X1 i_0_107 (.A(n_0_17), .B1(n_0_513), .B2(n_0_188), .ZN(n_0_125));
   AOI21_X1 i_0_108 (.A(n_0_483), .B1(n_0_198), .B2(n_0_127), .ZN(n_0_126));
   AOI221_X1 i_0_109 (.A(n_0_197), .B1(in_e[3]), .B2(in_m[15]), .C1(n_0_513), 
      .C2(in_m[7]), .ZN(n_0_127));
   AOI22_X1 i_0_110 (.A1(n_0_186), .A2(n_0_141), .B1(in_e[3]), .B2(n_0_20), 
      .ZN(n_0_128));
   NAND4_X1 i_0_111 (.A1(n_0_140), .A2(n_0_130), .A3(n_0_131), .A4(n_0_176), 
      .ZN(n_0_129));
   AOI22_X1 i_0_112 (.A1(n_0_13), .A2(n_0_310), .B1(in_e[2]), .B2(n_0_353), 
      .ZN(n_0_130));
   NAND2_X1 i_0_113 (.A1(n_0_14), .A2(n_0_322), .ZN(n_0_131));
   INV_X1 i_0_114 (.A(n_0_132), .ZN(n_4));
   AOI221_X1 i_0_115 (.A(n_0_167), .B1(n_0_162), .B2(n_0_133), .C1(in_e[4]), 
      .C2(n_0_136), .ZN(n_0_132));
   NAND2_X1 i_0_116 (.A1(n_0_135), .A2(n_0_134), .ZN(n_0_133));
   AOI22_X1 i_0_117 (.A1(n_0_33), .A2(n_0_160), .B1(n_0_32), .B2(n_0_156), 
      .ZN(n_0_134));
   AOI22_X1 i_0_118 (.A1(in_m[6]), .A2(n_0_30), .B1(n_0_31), .B2(n_0_433), 
      .ZN(n_0_135));
   NAND4_X1 i_0_119 (.A1(n_0_138), .A2(n_0_137), .A3(n_0_144), .A4(n_0_150), 
      .ZN(n_0_136));
   AOI21_X1 i_0_120 (.A(n_0_139), .B1(n_0_194), .B2(n_0_16), .ZN(n_0_137));
   NAND3_X1 i_0_121 (.A1(n_0_333), .A2(n_0_174), .A3(n_0_6), .ZN(n_0_138));
   NAND2_X1 i_0_122 (.A1(n_0_186), .A2(n_0_141), .ZN(n_0_16));
   NAND2_X1 i_0_123 (.A1(n_0_511), .A2(n_0_141), .ZN(n_0_17));
   AOI21_X1 i_0_124 (.A(n_0_142), .B1(n_0_141), .B2(n_0_140), .ZN(n_0_139));
   AOI22_X1 i_0_125 (.A1(n_0_12), .A2(n_0_309), .B1(n_0_351), .B2(n_0_19), 
      .ZN(n_0_140));
   INV_X1 i_0_126 (.A(n_0_18), .ZN(n_0_141));
   NAND2_X1 i_0_127 (.A1(n_0_513), .A2(n_0_512), .ZN(n_0_18));
   AOI21_X1 i_0_128 (.A(n_0_143), .B1(n_0_479), .B2(n_0_373), .ZN(n_0_142));
   AOI21_X1 i_0_129 (.A(n_0_308), .B1(n_0_513), .B2(n_0_487), .ZN(n_0_143));
   AOI221_X1 i_0_130 (.A(n_0_149), .B1(n_0_435), .B2(n_0_145), .C1(n_0_13), 
      .C2(n_0_310), .ZN(n_0_144));
   NAND3_X1 i_0_131 (.A1(n_0_147), .A2(n_0_146), .A3(n_0_148), .ZN(n_0_145));
   AOI222_X1 i_0_132 (.A1(n_0_5), .A2(n_0_296), .B1(n_0_4), .B2(n_0_315), 
      .C1(in_m[14]), .C2(n_0_2), .ZN(n_0_146));
   AOI22_X1 i_0_133 (.A1(n_0_3), .A2(n_0_347), .B1(n_0_0), .B2(n_0_383), 
      .ZN(n_0_147));
   NAND2_X1 i_0_134 (.A1(n_0_1), .A2(n_0_360), .ZN(n_0_148));
   AOI21_X1 i_0_135 (.A(n_0_513), .B1(n_0_311), .B2(n_0_263), .ZN(n_0_149));
   OAI22_X1 i_0_136 (.A1(n_0_404), .A2(n_0_322), .B1(in_e[3]), .B2(n_0_187), 
      .ZN(n_0_150));
   INV_X1 i_0_137 (.A(n_0_151), .ZN(n_5));
   AOI21_X1 i_0_138 (.A(n_0_153), .B1(in_e[5]), .B2(n_0_154), .ZN(n_0_151));
   OAI21_X1 i_0_139 (.A(n_0_152), .B1(n_0_514), .B2(n_0_153), .ZN(n_6));
   XNOR2_X1 i_0_140 (.A(in_e[7]), .B(n_0_152), .ZN(n_7));
   NAND2_X1 i_0_141 (.A1(n_0_514), .A2(n_0_153), .ZN(n_0_152));
   NOR2_X1 i_0_142 (.A1(in_e[5]), .A2(n_0_154), .ZN(n_0_153));
   AOI21_X1 i_0_143 (.A(n_0_167), .B1(n_0_162), .B2(n_0_155), .ZN(n_0_154));
   OAI221_X1 i_0_144 (.A(n_0_158), .B1(n_0_9), .B2(n_0_157), .C1(n_0_10), 
      .C2(n_0_161), .ZN(n_0_155));
   INV_X1 i_0_145 (.A(n_0_157), .ZN(n_0_156));
   NAND2_X1 i_0_146 (.A1(in_m[4]), .A2(n_0_393), .ZN(n_0_157));
   INV_X1 i_0_147 (.A(n_0_159), .ZN(n_0_158));
   OAI22_X1 i_0_148 (.A1(n_0_8), .A2(n_0_434), .B1(n_0_494), .B2(n_0_7), 
      .ZN(n_0_159));
   INV_X1 i_0_149 (.A(n_0_161), .ZN(n_0_160));
   NAND3_X1 i_0_150 (.A1(n_0_492), .A2(n_0_393), .A3(in_m[3]), .ZN(n_0_161));
   AND2_X1 i_0_151 (.A1(n_0_196), .A2(n_0_163), .ZN(n_0_162));
   AND2_X1 i_0_152 (.A1(n_0_329), .A2(n_0_164), .ZN(n_0_163));
   NOR2_X1 i_0_153 (.A1(in_m[12]), .A2(n_0_165), .ZN(n_0_164));
   NAND2_X1 i_0_154 (.A1(n_0_502), .A2(n_0_166), .ZN(n_0_165));
   NOR2_X1 i_0_155 (.A1(in_m[16]), .A2(n_0_324), .ZN(n_0_166));
   AOI21_X1 i_0_156 (.A(in_e[4]), .B1(n_0_177), .B2(n_0_168), .ZN(n_0_167));
   AND2_X1 i_0_157 (.A1(n_0_176), .A2(n_0_169), .ZN(n_0_168));
   AOI222_X1 i_0_158 (.A1(n_0_435), .A2(n_0_170), .B1(n_0_488), .B2(n_0_245), 
      .C1(n_0_174), .C2(n_0_173), .ZN(n_0_169));
   OAI221_X1 i_0_159 (.A(n_0_171), .B1(n_0_3), .B2(n_0_348), .C1(n_0_4), 
      .C2(n_0_316), .ZN(n_0_170));
   INV_X1 i_0_160 (.A(n_0_172), .ZN(n_0_171));
   OAI22_X1 i_0_161 (.A1(n_0_0), .A2(n_0_384), .B1(n_0_1), .B2(n_0_361), 
      .ZN(n_0_172));
   OAI22_X1 i_0_162 (.A1(n_0_6), .A2(n_0_334), .B1(n_0_5), .B2(n_0_423), 
      .ZN(n_0_173));
   INV_X1 i_0_163 (.A(n_0_175), .ZN(n_0_174));
   NAND2_X1 i_0_164 (.A1(n_0_451), .A2(n_0_435), .ZN(n_0_175));
   NAND2_X1 i_0_165 (.A1(n_0_451), .A2(n_0_327), .ZN(n_0_176));
   INV_X1 i_0_166 (.A(n_0_178), .ZN(n_0_177));
   AOI21_X1 i_0_167 (.A(in_e[3]), .B1(n_0_187), .B2(n_0_180), .ZN(n_0_178));
   AOI21_X1 i_0_168 (.A(n_0_182), .B1(n_0_485), .B2(n_0_322), .ZN(n_0_179));
   AOI221_X1 i_0_169 (.A(n_0_182), .B1(n_0_351), .B2(n_0_181), .C1(n_0_194), 
      .C2(n_0_185), .ZN(n_0_180));
   INV_X1 i_0_170 (.A(n_0_181), .ZN(n_0_19));
   NOR2_X1 i_0_171 (.A1(in_e[2]), .A2(n_0_11), .ZN(n_0_181));
   OAI211_X1 i_0_172 (.A(n_0_183), .B(n_0_184), .C1(n_0_13), .C2(n_0_311), 
      .ZN(n_0_182));
   NAND2_X1 i_0_173 (.A1(n_0_512), .A2(n_0_353), .ZN(n_0_183));
   AOI21_X1 i_0_174 (.A(n_0_264), .B1(n_0_487), .B2(n_0_309), .ZN(n_0_184));
   INV_X1 i_0_175 (.A(n_0_20), .ZN(n_0_185));
   NAND2_X1 i_0_176 (.A1(n_0_510), .A2(n_0_188), .ZN(n_0_20));
   INV_X1 i_0_177 (.A(n_0_21), .ZN(n_0_186));
   NAND2_X1 i_0_178 (.A1(n_0_511), .A2(n_0_510), .ZN(n_0_21));
   AOI22_X1 i_0_179 (.A1(n_0_485), .A2(n_0_322), .B1(n_0_404), .B2(n_0_188), 
      .ZN(n_0_187));
   INV_X1 i_0_180 (.A(n_0_22), .ZN(n_0_188));
   NAND2_X1 i_0_181 (.A1(n_0_512), .A2(n_0_511), .ZN(n_0_22));
   AOI21_X1 i_0_182 (.A(in_m[23]), .B1(n_0_340), .B2(n_0_189), .ZN(n_8));
   NOR4_X1 i_0_183 (.A1(in_m[22]), .A2(in_m[15]), .A3(n_0_190), .A4(n_0_191), 
      .ZN(n_0_189));
   NAND3_X1 i_0_184 (.A1(n_0_509), .A2(n_0_475), .A3(n_0_393), .ZN(n_0_190));
   NAND4_X1 i_0_185 (.A1(n_0_492), .A2(n_0_491), .A3(n_0_498), .A4(n_0_201), 
      .ZN(n_0_191));
   AND2_X1 i_0_186 (.A1(in_m[0]), .A2(n_0_194), .ZN(n_9));
   OAI21_X1 i_0_187 (.A(n_0_192), .B1(n_0_489), .B2(n_0_195), .ZN(n_10));
   NAND2_X1 i_0_188 (.A1(in_m[0]), .A2(n_0_404), .ZN(n_0_192));
   OAI21_X1 i_0_189 (.A(n_0_193), .B1(n_0_490), .B2(n_0_195), .ZN(n_11));
   AOI22_X1 i_0_190 (.A1(in_m[0]), .A2(n_0_351), .B1(in_m[1]), .B2(n_0_404), 
      .ZN(n_0_193));
   INV_X1 i_0_191 (.A(n_0_195), .ZN(n_0_194));
   AOI21_X1 i_0_192 (.A(n_0_483), .B1(n_0_198), .B2(n_0_196), .ZN(n_0_195));
   NOR3_X1 i_0_193 (.A1(in_m[15]), .A2(in_m[7]), .A3(n_0_197), .ZN(n_0_196));
   NAND4_X1 i_0_194 (.A1(n_0_501), .A2(n_0_499), .A3(n_0_509), .A4(n_0_475), 
      .ZN(n_0_197));
   NOR2_X1 i_0_195 (.A1(in_m[3]), .A2(n_0_199), .ZN(n_0_198));
   NAND3_X1 i_0_196 (.A1(n_0_466), .A2(n_0_201), .A3(n_0_200), .ZN(n_0_199));
   NOR3_X1 i_0_197 (.A1(in_m[4]), .A2(n_0_394), .A3(n_0_330), .ZN(n_0_200));
   NOR3_X1 i_0_198 (.A1(in_m[20]), .A2(in_m[18]), .A3(in_m[16]), .ZN(n_0_201));
   OAI221_X1 i_0_199 (.A(n_0_202), .B1(n_0_490), .B2(n_0_405), .C1(n_0_491), 
      .C2(n_0_484), .ZN(n_12));
   AOI22_X1 i_0_200 (.A1(in_m[0]), .A2(n_0_353), .B1(in_m[1]), .B2(n_0_351), 
      .ZN(n_0_202));
   OAI211_X1 i_0_201 (.A(n_0_204), .B(n_0_203), .C1(n_0_492), .C2(n_0_484), 
      .ZN(n_13));
   AOI22_X1 i_0_202 (.A1(in_m[0]), .A2(n_0_309), .B1(in_m[2]), .B2(n_0_351), 
      .ZN(n_0_203));
   AOI22_X1 i_0_203 (.A1(in_m[1]), .A2(n_0_353), .B1(in_m[3]), .B2(n_0_404), 
      .ZN(n_0_204));
   OAI211_X1 i_0_204 (.A(n_0_206), .B(n_0_205), .C1(n_0_492), .C2(n_0_405), 
      .ZN(n_14));
   AOI222_X1 i_0_205 (.A1(in_m[3]), .A2(n_0_351), .B1(in_m[5]), .B2(n_0_483), 
      .C1(in_m[2]), .C2(n_0_353), .ZN(n_0_205));
   AOI22_X1 i_0_206 (.A1(in_m[0]), .A2(n_0_310), .B1(in_m[1]), .B2(n_0_309), 
      .ZN(n_0_206));
   NAND2_X1 i_0_207 (.A1(n_0_209), .A2(n_0_207), .ZN(n_15));
   AOI221_X1 i_0_208 (.A(n_0_208), .B1(in_m[1]), .B2(n_0_310), .C1(in_m[0]), 
      .C2(n_0_322), .ZN(n_0_207));
   OAI222_X1 i_0_209 (.A1(n_0_493), .A2(n_0_405), .B1(n_0_494), .B2(n_0_484), 
      .C1(n_0_492), .C2(n_0_352), .ZN(n_0_208));
   AOI22_X1 i_0_210 (.A1(in_m[2]), .A2(n_0_309), .B1(in_m[3]), .B2(n_0_353), 
      .ZN(n_0_209));
   NAND3_X1 i_0_211 (.A1(n_0_211), .A2(n_0_210), .A3(n_0_212), .ZN(n_16));
   AOI22_X1 i_0_212 (.A1(in_m[1]), .A2(n_0_322), .B1(in_m[4]), .B2(n_0_353), 
      .ZN(n_0_210));
   AOI222_X1 i_0_213 (.A1(in_m[0]), .A2(n_0_264), .B1(in_m[7]), .B2(n_0_483), 
      .C1(in_m[5]), .C2(n_0_351), .ZN(n_0_211));
   AOI222_X1 i_0_214 (.A1(in_m[2]), .A2(n_0_310), .B1(in_m[3]), .B2(n_0_309), 
      .C1(in_m[6]), .C2(n_0_404), .ZN(n_0_212));
   OAI221_X1 i_0_215 (.A(n_0_213), .B1(n_0_491), .B2(n_0_311), .C1(n_0_490), 
      .C2(n_0_323), .ZN(n_17));
   AOI221_X1 i_0_216 (.A(n_0_214), .B1(in_m[4]), .B2(n_0_309), .C1(in_m[6]), 
      .C2(n_0_351), .ZN(n_0_213));
   OAI221_X1 i_0_217 (.A(n_0_215), .B1(n_0_502), .B2(n_0_321), .C1(n_0_489), 
      .C2(n_0_263), .ZN(n_0_214));
   AOI222_X1 i_0_218 (.A1(in_m[7]), .A2(n_0_404), .B1(in_m[5]), .B2(n_0_353), 
      .C1(in_m[8]), .C2(n_0_483), .ZN(n_0_215));
   NAND4_X1 i_0_219 (.A1(n_0_219), .A2(n_0_216), .A3(n_0_218), .A4(n_0_217), 
      .ZN(n_18));
   AOI222_X1 i_0_220 (.A1(in_m[2]), .A2(n_0_264), .B1(in_m[0]), .B2(n_0_240), 
      .C1(in_m[1]), .C2(n_0_245), .ZN(n_0_216));
   AOI22_X1 i_0_221 (.A1(in_m[4]), .A2(n_0_310), .B1(in_m[3]), .B2(n_0_322), 
      .ZN(n_0_217));
   AOI22_X1 i_0_222 (.A1(in_m[6]), .A2(n_0_353), .B1(in_m[5]), .B2(n_0_309), 
      .ZN(n_0_218));
   AOI222_X1 i_0_223 (.A1(in_m[9]), .A2(n_0_483), .B1(in_m[8]), .B2(n_0_404), 
      .C1(in_m[7]), .C2(n_0_351), .ZN(n_0_219));
   OAI211_X1 i_0_224 (.A(n_0_220), .B(n_0_221), .C1(n_0_492), .C2(n_0_323), 
      .ZN(n_19));
   AOI222_X1 i_0_225 (.A1(in_m[1]), .A2(n_0_240), .B1(in_m[2]), .B2(n_0_245), 
      .C1(n_0_383), .C2(n_0_320), .ZN(n_0_220));
   AOI21_X1 i_0_226 (.A(n_0_222), .B1(in_m[3]), .B2(n_0_264), .ZN(n_0_221));
   OAI211_X1 i_0_227 (.A(n_0_223), .B(n_0_224), .C1(n_0_493), .C2(n_0_311), 
      .ZN(n_0_222));
   AOI222_X1 i_0_228 (.A1(in_m[10]), .A2(n_0_483), .B1(in_m[9]), .B2(n_0_404), 
      .C1(in_m[8]), .C2(n_0_351), .ZN(n_0_223));
   AOI22_X1 i_0_229 (.A1(in_m[7]), .A2(n_0_353), .B1(in_m[6]), .B2(n_0_309), 
      .ZN(n_0_224));
   OAI211_X1 i_0_230 (.A(n_0_225), .B(n_0_229), .C1(n_0_495), .C2(n_0_308), 
      .ZN(n_20));
   AOI221_X1 i_0_231 (.A(n_0_228), .B1(n_0_435), .B2(n_0_227), .C1(in_m[0]), 
      .C2(n_0_226), .ZN(n_0_225));
   NOR2_X1 i_0_232 (.A1(n_0_348), .A2(n_0_260), .ZN(n_0_226));
   OAI222_X1 i_0_233 (.A1(n_0_502), .A2(n_0_491), .B1(n_0_490), .B2(n_0_361), 
      .C1(n_0_489), .C2(n_0_384), .ZN(n_0_227));
   OAI221_X1 i_0_234 (.A(n_0_230), .B1(n_0_497), .B2(n_0_352), .C1(n_0_492), 
      .C2(n_0_263), .ZN(n_0_228));
   AOI222_X1 i_0_235 (.A1(in_m[6]), .A2(n_0_310), .B1(in_m[8]), .B2(n_0_353), 
      .C1(in_m[5]), .C2(n_0_322), .ZN(n_0_229));
   AOI22_X1 i_0_236 (.A1(in_m[10]), .A2(n_0_404), .B1(in_m[11]), .B2(n_0_483), 
      .ZN(n_0_230));
   NAND4_X1 i_0_237 (.A1(n_0_235), .A2(n_0_231), .A3(n_0_237), .A4(n_0_238), 
      .ZN(n_21));
   INV_X1 i_0_238 (.A(n_0_232), .ZN(n_0_231));
   OAI211_X1 i_0_239 (.A(n_0_234), .B(n_0_233), .C1(n_0_500), .C2(n_0_484), 
      .ZN(n_0_232));
   AOI22_X1 i_0_240 (.A1(in_m[5]), .A2(n_0_264), .B1(in_m[4]), .B2(n_0_245), 
      .ZN(n_0_233));
   AOI22_X1 i_0_241 (.A1(in_m[11]), .A2(n_0_404), .B1(in_m[9]), .B2(n_0_353), 
      .ZN(n_0_234));
   AOI221_X1 i_0_242 (.A(n_0_236), .B1(in_m[7]), .B2(n_0_310), .C1(in_m[8]), 
      .C2(n_0_309), .ZN(n_0_235));
   OAI33_X1 i_0_243 (.A1(n_0_348), .A2(n_0_257), .A3(n_0_489), .B1(n_0_384), 
      .B2(n_0_260), .B3(n_0_490), .ZN(n_0_236));
   NAND2_X1 i_0_244 (.A1(in_m[6]), .A2(n_0_322), .ZN(n_0_237));
   AOI22_X1 i_0_245 (.A1(in_m[3]), .A2(n_0_240), .B1(in_m[10]), .B2(n_0_239), 
      .ZN(n_0_238));
   OAI21_X1 i_0_246 (.A(n_0_352), .B1(n_0_379), .B2(n_0_332), .ZN(n_0_239));
   NOR2_X1 i_0_247 (.A1(n_0_436), .A2(n_0_361), .ZN(n_0_240));
   NAND4_X1 i_0_248 (.A1(n_0_246), .A2(n_0_244), .A3(n_0_243), .A4(n_0_241), 
      .ZN(n_22));
   AOI21_X1 i_0_249 (.A(n_0_242), .B1(in_m[6]), .B2(n_0_264), .ZN(n_0_241));
   NOR3_X1 i_0_250 (.A1(n_0_489), .A2(n_0_316), .A3(n_0_290), .ZN(n_0_242));
   NAND4_X1 i_0_251 (.A1(n_0_475), .A2(n_0_438), .A3(in_m[0]), .A4(n_0_296), 
      .ZN(n_0_243));
   AOI22_X1 i_0_252 (.A1(in_m[7]), .A2(n_0_322), .B1(in_m[5]), .B2(n_0_245), 
      .ZN(n_0_244));
   NOR2_X1 i_0_253 (.A1(n_0_502), .A2(n_0_436), .ZN(n_0_245));
   AOI211_X1 i_0_254 (.A(n_0_251), .B(n_0_247), .C1(in_m[9]), .C2(n_0_309), 
      .ZN(n_0_246));
   OAI211_X1 i_0_255 (.A(n_0_250), .B(n_0_248), .C1(n_0_496), .C2(n_0_311), 
      .ZN(n_0_247));
   AOI21_X1 i_0_256 (.A(n_0_249), .B1(in_m[10]), .B2(n_0_353), .ZN(n_0_248));
   NOR3_X1 i_0_257 (.A1(n_0_491), .A2(n_0_384), .A3(n_0_257), .ZN(n_0_249));
   AOI222_X1 i_0_258 (.A1(in_m[13]), .A2(n_0_483), .B1(in_m[12]), .B2(n_0_404), 
      .C1(in_m[11]), .C2(n_0_351), .ZN(n_0_250));
   OAI33_X1 i_0_259 (.A1(n_0_492), .A2(n_0_361), .A3(n_0_260), .B1(n_0_490), 
      .B2(n_0_348), .B3(n_0_379), .ZN(n_0_251));
   NAND4_X1 i_0_260 (.A1(n_0_255), .A2(n_0_252), .A3(n_0_258), .A4(n_0_261), 
      .ZN(n_23));
   AOI211_X1 i_0_261 (.A(n_0_253), .B(n_0_254), .C1(in_m[10]), .C2(n_0_309), 
      .ZN(n_0_252));
   OAI22_X1 i_0_262 (.A1(n_0_500), .A2(n_0_352), .B1(n_0_501), .B2(n_0_405), 
      .ZN(n_0_253));
   NOR3_X1 i_0_263 (.A1(n_0_334), .A2(n_0_332), .A3(n_0_411), .ZN(n_0_254));
   AOI221_X1 i_0_264 (.A(n_0_256), .B1(in_m[11]), .B2(n_0_353), .C1(in_m[9]), 
      .C2(n_0_310), .ZN(n_0_255));
   OAI33_X1 i_0_265 (.A1(n_0_493), .A2(n_0_361), .A3(n_0_257), .B1(n_0_492), 
      .B2(n_0_384), .B3(n_0_379), .ZN(n_0_256));
   NAND2_X1 i_0_266 (.A1(n_0_481), .A2(n_0_437), .ZN(n_0_257));
   AOI22_X1 i_0_267 (.A1(in_m[8]), .A2(n_0_322), .B1(in_m[14]), .B2(n_0_259), 
      .ZN(n_0_258));
   OAI21_X1 i_0_268 (.A(n_0_484), .B1(n_0_494), .B2(n_0_260), .ZN(n_0_259));
   NAND2_X1 i_0_269 (.A1(n_0_437), .A2(n_0_356), .ZN(n_0_260));
   AOI211_X1 i_0_270 (.A(n_0_265), .B(n_0_262), .C1(in_m[7]), .C2(n_0_264), 
      .ZN(n_0_261));
   OAI33_X1 i_0_271 (.A1(n_0_489), .A2(n_0_297), .A3(n_0_377), .B1(n_0_490), 
      .B2(n_0_316), .B3(n_0_357), .ZN(n_0_262));
   INV_X1 i_0_272 (.A(n_0_264), .ZN(n_0_263));
   NOR2_X1 i_0_273 (.A1(n_0_483), .A2(n_0_278), .ZN(n_0_264));
   NOR3_X1 i_0_274 (.A1(n_0_491), .A2(n_0_348), .A3(n_0_290), .ZN(n_0_265));
   NAND4_X1 i_0_275 (.A1(n_0_272), .A2(n_0_271), .A3(n_0_275), .A4(n_0_266), 
      .ZN(n_24));
   AOI211_X1 i_0_276 (.A(n_0_267), .B(n_0_268), .C1(in_m[9]), .C2(n_0_322), 
      .ZN(n_0_266));
   NOR3_X1 i_0_277 (.A1(n_0_384), .A2(n_0_290), .A3(n_0_493), .ZN(n_0_267));
   OAI211_X1 i_0_278 (.A(n_0_269), .B(n_0_270), .C1(n_0_379), .C2(n_0_280), 
      .ZN(n_0_268));
   AOI22_X1 i_0_279 (.A1(in_m[12]), .A2(n_0_353), .B1(in_m[11]), .B2(n_0_309), 
      .ZN(n_0_269));
   AOI222_X1 i_0_280 (.A1(in_m[13]), .A2(n_0_351), .B1(in_m[10]), .B2(n_0_310), 
      .C1(in_m[15]), .C2(n_0_483), .ZN(n_0_270));
   NAND4_X1 i_0_281 (.A1(n_0_501), .A2(n_0_453), .A3(n_0_327), .A4(in_m[0]), 
      .ZN(n_0_271));
   NOR3_X1 i_0_282 (.A1(n_0_279), .A2(n_0_273), .A3(n_0_274), .ZN(n_0_272));
   NOR3_X1 i_0_283 (.A1(n_0_357), .A2(n_0_348), .A3(n_0_492), .ZN(n_0_273));
   OAI33_X1 i_0_284 (.A1(n_0_490), .A2(n_0_297), .A3(n_0_411), .B1(n_0_491), 
      .B2(n_0_377), .B3(n_0_316), .ZN(n_0_274));
   INV_X1 i_0_285 (.A(n_0_276), .ZN(n_0_275));
   AOI21_X1 i_0_286 (.A(n_0_496), .B1(n_0_278), .B2(n_0_277), .ZN(n_0_276));
   NAND4_X1 i_0_287 (.A1(in_m[1]), .A2(n_0_415), .A3(n_0_447), .A4(n_0_451), 
      .ZN(n_0_277));
   NAND3_X1 i_0_288 (.A1(n_0_504), .A2(in_m[15]), .A3(n_0_293), .ZN(n_0_278));
   AOI21_X1 i_0_289 (.A(n_0_502), .B1(n_0_405), .B2(n_0_364), .ZN(n_0_279));
   NAND2_X1 i_0_290 (.A1(in_m[6]), .A2(n_0_360), .ZN(n_0_280));
   OR3_X1 i_0_291 (.A1(n_0_295), .A2(n_0_281), .A3(n_0_288), .ZN(n_25));
   NAND2_X1 i_0_292 (.A1(n_0_286), .A2(n_0_282), .ZN(n_0_281));
   AOI211_X1 i_0_293 (.A(n_0_285), .B(n_0_283), .C1(in_m[15]), .C2(n_0_300), 
      .ZN(n_0_282));
   OAI211_X1 i_0_294 (.A(n_0_294), .B(n_0_284), .C1(n_0_500), .C2(n_0_308), 
      .ZN(n_0_283));
   AOI21_X1 i_0_295 (.A(n_0_289), .B1(in_m[11]), .B2(n_0_310), .ZN(n_0_284));
   OAI33_X1 i_0_296 (.A1(n_0_321), .A2(n_0_298), .A3(n_0_494), .B1(n_0_411), 
      .B2(n_0_316), .B3(n_0_492), .ZN(n_0_285));
   AOI211_X1 i_0_297 (.A(n_0_287), .B(n_0_299), .C1(in_m[16]), .C2(n_0_291), 
      .ZN(n_0_286));
   OAI33_X1 i_0_298 (.A1(n_0_361), .A2(n_0_290), .A3(n_0_495), .B1(n_0_384), 
      .B2(n_0_357), .B3(n_0_494), .ZN(n_0_287));
   OAI33_X1 i_0_299 (.A1(n_0_416), .A2(n_0_297), .A3(n_0_491), .B1(n_0_362), 
      .B2(n_0_330), .B3(n_0_489), .ZN(n_0_288));
   NOR4_X1 i_0_300 (.A1(n_0_338), .A2(n_0_334), .A3(n_0_490), .A4(n_0_436), 
      .ZN(n_0_289));
   NAND2_X1 i_0_301 (.A1(n_0_438), .A2(n_0_370), .ZN(n_0_290));
   INV_X1 i_0_302 (.A(n_0_292), .ZN(n_0_291));
   AOI21_X1 i_0_303 (.A(n_0_483), .B1(in_m[10]), .B2(n_0_293), .ZN(n_0_292));
   AND2_X1 i_0_304 (.A1(n_0_473), .A2(n_0_356), .ZN(n_0_293));
   NAND2_X1 i_0_305 (.A1(in_m[13]), .A2(n_0_353), .ZN(n_0_294));
   AOI21_X1 i_0_306 (.A(n_0_502), .B1(n_0_378), .B2(n_0_352), .ZN(n_0_295));
   INV_X1 i_0_307 (.A(n_0_297), .ZN(n_0_296));
   NAND2_X1 i_0_308 (.A1(n_0_451), .A2(n_0_422), .ZN(n_0_297));
   NAND3_X1 i_0_309 (.A1(n_0_426), .A2(n_0_329), .A3(n_0_495), .ZN(n_0_298));
   NOR3_X1 i_0_310 (.A1(n_0_493), .A2(n_0_348), .A3(n_0_377), .ZN(n_0_299));
   OAI21_X1 i_0_311 (.A(n_0_405), .B1(n_0_497), .B2(n_0_416), .ZN(n_0_300));
   NAND3_X1 i_0_312 (.A1(n_0_306), .A2(n_0_301), .A3(n_0_317), .ZN(n_26));
   NOR4_X1 i_0_313 (.A1(n_0_305), .A2(n_0_304), .A3(n_0_325), .A4(n_0_302), 
      .ZN(n_0_301));
   AOI21_X1 i_0_314 (.A(n_0_436), .B1(n_0_312), .B2(n_0_303), .ZN(n_0_302));
   NAND3_X1 i_0_315 (.A1(in_m[0]), .A2(n_0_340), .A3(n_0_433), .ZN(n_0_303));
   OAI222_X1 i_0_316 (.A1(n_0_499), .A2(n_0_323), .B1(n_0_504), .B2(n_0_405), 
      .C1(n_0_505), .C2(n_0_484), .ZN(n_0_304));
   OAI33_X1 i_0_317 (.A1(n_0_411), .A2(n_0_348), .A3(n_0_494), .B1(n_0_416), 
      .B2(n_0_316), .B3(n_0_493), .ZN(n_0_305));
   AOI221_X1 i_0_318 (.A(n_0_307), .B1(in_m[12]), .B2(n_0_310), .C1(in_m[13]), 
      .C2(n_0_309), .ZN(n_0_306));
   OAI33_X1 i_0_319 (.A1(n_0_384), .A2(n_0_377), .A3(n_0_495), .B1(n_0_361), 
      .B2(n_0_357), .B3(n_0_496), .ZN(n_0_307));
   INV_X1 i_0_320 (.A(n_0_309), .ZN(n_0_308));
   NOR2_X1 i_0_321 (.A1(n_0_483), .A2(n_0_355), .ZN(n_0_309));
   INV_X1 i_0_322 (.A(n_0_311), .ZN(n_0_310));
   NAND3_X1 i_0_323 (.A1(in_m[17]), .A2(n_0_477), .A3(n_0_474), .ZN(n_0_311));
   AOI21_X1 i_0_324 (.A(n_0_313), .B1(n_0_329), .B2(n_0_314), .ZN(n_0_312));
   OAI33_X1 i_0_325 (.A1(n_0_363), .A2(n_0_334), .A3(n_0_491), .B1(n_0_423), 
      .B2(n_0_338), .B3(n_0_492), .ZN(n_0_313));
   NOR4_X1 i_0_326 (.A1(n_0_489), .A2(n_0_425), .A3(in_m[7]), .A4(n_0_494), 
      .ZN(n_0_314));
   INV_X1 i_0_327 (.A(n_0_316), .ZN(n_0_315));
   NAND2_X1 i_0_328 (.A1(in_m[10]), .A2(n_0_451), .ZN(n_0_316));
   AOI22_X1 i_0_329 (.A1(in_m[14]), .A2(n_0_319), .B1(in_m[15]), .B2(n_0_318), 
      .ZN(n_0_317));
   OAI21_X1 i_0_330 (.A(n_0_352), .B1(n_0_498), .B2(n_0_416), .ZN(n_0_318));
   OAI22_X1 i_0_331 (.A1(n_0_497), .A2(n_0_436), .B1(n_0_507), .B2(n_0_478), 
      .ZN(n_0_319));
   INV_X1 i_0_332 (.A(n_0_321), .ZN(n_0_320));
   NAND2_X1 i_0_333 (.A1(in_m[0]), .A2(n_0_435), .ZN(n_0_321));
   INV_X1 i_0_334 (.A(n_0_323), .ZN(n_0_322));
   NAND3_X1 i_0_335 (.A1(n_0_506), .A2(n_0_481), .A3(n_0_412), .ZN(n_0_323));
   NAND2_X1 i_0_336 (.A1(n_0_506), .A2(n_0_481), .ZN(n_0_324));
   NOR4_X1 i_0_337 (.A1(n_0_427), .A2(n_0_330), .A3(n_0_490), .A4(n_0_364), 
      .ZN(n_0_325));
   OAI221_X1 i_0_338 (.A(n_0_341), .B1(n_0_491), .B2(n_0_326), .C1(n_0_436), 
      .C2(n_0_328), .ZN(n_27));
   NAND2_X1 i_0_339 (.A1(n_0_424), .A2(n_0_327), .ZN(n_0_326));
   NOR2_X1 i_0_340 (.A1(n_0_364), .A2(n_0_330), .ZN(n_0_327));
   AOI221_X1 i_0_341 (.A(n_0_331), .B1(n_0_498), .B2(n_0_335), .C1(in_m[6]), 
      .C2(n_0_337), .ZN(n_0_328));
   INV_X1 i_0_342 (.A(n_0_330), .ZN(n_0_329));
   NAND2_X1 i_0_343 (.A1(n_0_496), .A2(n_0_447), .ZN(n_0_330));
   OAI33_X1 i_0_344 (.A1(n_0_492), .A2(n_0_427), .A3(n_0_334), .B1(n_0_430), 
      .B2(n_0_394), .B3(n_0_332), .ZN(n_0_331));
   NAND2_X1 i_0_345 (.A1(in_m[0]), .A2(n_0_451), .ZN(n_0_332));
   INV_X1 i_0_346 (.A(n_0_334), .ZN(n_0_333));
   NAND2_X1 i_0_347 (.A1(in_m[8]), .A2(n_0_447), .ZN(n_0_334));
   AND2_X1 i_0_348 (.A1(in_m[5]), .A2(n_0_336), .ZN(n_0_335));
   OAI33_X1 i_0_349 (.A1(n_0_489), .A2(n_0_459), .A3(n_0_450), .B1(in_m[11]), 
      .B2(n_0_467), .B3(n_0_497), .ZN(n_0_336));
   OAI21_X1 i_0_350 (.A(n_0_339), .B1(n_0_498), .B2(n_0_338), .ZN(n_0_337));
   NAND2_X1 i_0_351 (.A1(n_0_501), .A2(n_0_453), .ZN(n_0_338));
   NAND2_X1 i_0_352 (.A1(in_m[2]), .A2(n_0_340), .ZN(n_0_339));
   NOR3_X1 i_0_353 (.A1(in_m[9]), .A2(in_m[7]), .A3(n_0_450), .ZN(n_0_340));
   AND4_X1 i_0_354 (.A1(n_0_344), .A2(n_0_342), .A3(n_0_345), .A4(n_0_346), 
      .ZN(n_0_341));
   INV_X1 i_0_355 (.A(n_0_343), .ZN(n_0_342));
   OAI33_X1 i_0_356 (.A1(n_0_416), .A2(n_0_348), .A3(n_0_495), .B1(n_0_377), 
      .B2(n_0_361), .B3(n_0_497), .ZN(n_0_343));
   AOI222_X1 i_0_357 (.A1(in_m[15]), .A2(n_0_353), .B1(in_m[18]), .B2(n_0_483), 
      .C1(n_0_370), .C2(n_0_350), .ZN(n_0_344));
   NAND3_X1 i_0_358 (.A1(in_m[8]), .A2(n_0_410), .A3(n_0_383), .ZN(n_0_345));
   AOI221_X1 i_0_359 (.A(n_0_349), .B1(in_m[14]), .B2(n_0_354), .C1(in_m[16]), 
      .C2(n_0_351), .ZN(n_0_346));
   INV_X1 i_0_360 (.A(n_0_348), .ZN(n_0_347));
   NAND2_X1 i_0_361 (.A1(in_m[11]), .A2(n_0_424), .ZN(n_0_348));
   AOI21_X1 i_0_362 (.A(n_0_505), .B1(n_0_407), .B2(n_0_405), .ZN(n_0_349));
   OAI33_X1 i_0_363 (.A1(n_0_499), .A2(n_0_408), .A3(n_0_478), .B1(n_0_500), 
      .B2(n_0_480), .B3(n_0_442), .ZN(n_0_350));
   INV_X1 i_0_364 (.A(n_0_352), .ZN(n_0_351));
   NAND2_X1 i_0_365 (.A1(in_m[20]), .A2(n_0_479), .ZN(n_0_352));
   NOR2_X1 i_0_366 (.A1(n_0_507), .A2(n_0_478), .ZN(n_0_353));
   OAI21_X1 i_0_367 (.A(n_0_355), .B1(n_0_498), .B2(n_0_357), .ZN(n_0_354));
   NAND2_X1 i_0_368 (.A1(in_m[18]), .A2(n_0_356), .ZN(n_0_355));
   NOR2_X1 i_0_369 (.A1(in_m[21]), .A2(n_0_373), .ZN(n_0_356));
   NAND2_X1 i_0_370 (.A1(n_0_475), .A2(n_0_438), .ZN(n_0_357));
   NAND4_X1 i_0_371 (.A1(n_0_380), .A2(n_0_374), .A3(n_0_365), .A4(n_0_358), 
      .ZN(n_28));
   AOI22_X1 i_0_372 (.A1(n_0_479), .A2(n_0_366), .B1(in_m[10]), .B2(n_0_359), 
      .ZN(n_0_358));
   OAI21_X1 i_0_373 (.A(n_0_362), .B1(n_0_411), .B2(n_0_361), .ZN(n_0_359));
   INV_X1 i_0_374 (.A(n_0_361), .ZN(n_0_360));
   NAND2_X1 i_0_375 (.A1(n_0_502), .A2(in_m[13]), .ZN(n_0_361));
   OR2_X1 i_0_376 (.A1(n_0_364), .A2(n_0_363), .ZN(n_0_362));
   NAND2_X1 i_0_377 (.A1(n_0_499), .A2(n_0_466), .ZN(n_0_363));
   NAND2_X1 i_0_378 (.A1(in_m[7]), .A2(n_0_435), .ZN(n_0_364));
   NAND3_X1 i_0_379 (.A1(in_m[18]), .A2(n_0_484), .A3(n_0_372), .ZN(n_0_365));
   OAI21_X1 i_0_380 (.A(n_0_368), .B1(n_0_505), .B2(n_0_367), .ZN(n_0_366));
   AOI21_X1 i_0_381 (.A(in_m[20]), .B1(in_m[14]), .B2(n_0_474), .ZN(n_0_367));
   NAND2_X1 i_0_382 (.A1(n_0_508), .A2(n_0_369), .ZN(n_0_368));
   OAI33_X1 i_0_383 (.A1(n_0_476), .A2(n_0_408), .A3(n_0_500), .B1(n_0_501), 
      .B2(n_0_371), .B3(n_0_504), .ZN(n_0_369));
   INV_X1 i_0_384 (.A(n_0_371), .ZN(n_0_370));
   NAND2_X1 i_0_385 (.A1(n_0_506), .A2(n_0_505), .ZN(n_0_371));
   OAI21_X1 i_0_386 (.A(n_0_509), .B1(n_0_503), .B2(n_0_373), .ZN(n_0_372));
   NAND2_X1 i_0_387 (.A1(n_0_508), .A2(n_0_507), .ZN(n_0_373));
   OAI21_X1 i_0_388 (.A(in_m[11]), .B1(n_0_376), .B2(n_0_375), .ZN(n_0_374));
   NOR4_X1 i_0_389 (.A1(in_m[20]), .A2(n_0_378), .A3(in_m[12]), .A4(in_m[13]), 
      .ZN(n_0_375));
   NOR2_X1 i_0_390 (.A1(n_0_502), .A2(n_0_377), .ZN(n_0_376));
   NAND2_X1 i_0_391 (.A1(n_0_474), .A2(n_0_438), .ZN(n_0_377));
   NAND3_X1 i_0_392 (.A1(n_0_479), .A2(n_0_437), .A3(in_m[8]), .ZN(n_0_378));
   NAND2_X1 i_0_393 (.A1(n_0_479), .A2(n_0_437), .ZN(n_0_379));
   AOI221_X1 i_0_394 (.A(n_0_382), .B1(in_m[19]), .B2(n_0_381), .C1(n_0_435), 
      .C2(n_0_385), .ZN(n_0_380));
   OAI21_X1 i_0_395 (.A(n_0_484), .B1(n_0_504), .B2(n_0_478), .ZN(n_0_381));
   NOR3_X1 i_0_396 (.A1(n_0_497), .A2(n_0_416), .A3(n_0_384), .ZN(n_0_382));
   INV_X1 i_0_397 (.A(n_0_384), .ZN(n_0_383));
   NAND2_X1 i_0_398 (.A1(in_m[12]), .A2(n_0_454), .ZN(n_0_384));
   OAI211_X1 i_0_399 (.A(n_0_389), .B(n_0_386), .C1(n_0_450), .C2(n_0_390), 
      .ZN(n_0_385));
   NAND3_X1 i_0_400 (.A1(n_0_447), .A2(n_0_424), .A3(n_0_387), .ZN(n_0_386));
   AOI21_X1 i_0_401 (.A(n_0_493), .B1(n_0_496), .B2(n_0_388), .ZN(n_0_387));
   NAND3_X1 i_0_402 (.A1(n_0_499), .A2(in_m[2]), .A3(n_0_458), .ZN(n_0_388));
   NAND3_X1 i_0_403 (.A1(in_m[6]), .A2(n_0_422), .A3(n_0_426), .ZN(n_0_389));
   AOI22_X1 i_0_404 (.A1(n_0_498), .A2(n_0_395), .B1(n_0_497), .B2(n_0_391), 
      .ZN(n_0_390));
   AOI21_X1 i_0_405 (.A(n_0_492), .B1(n_0_495), .B2(n_0_392), .ZN(n_0_391));
   NAND3_X1 i_0_406 (.A1(n_0_498), .A2(in_m[1]), .A3(n_0_393), .ZN(n_0_392));
   INV_X1 i_0_407 (.A(n_0_394), .ZN(n_0_393));
   NAND2_X1 i_0_408 (.A1(n_0_494), .A2(n_0_493), .ZN(n_0_394));
   AOI211_X1 i_0_409 (.A(in_m[7]), .B(n_0_491), .C1(n_0_494), .C2(n_0_396), 
      .ZN(n_0_395));
   NAND4_X1 i_0_410 (.A1(n_0_497), .A2(n_0_493), .A3(n_0_492), .A4(in_m[0]), 
      .ZN(n_0_396));
   OAI211_X1 i_0_411 (.A(n_0_413), .B(n_0_397), .C1(n_0_436), .C2(n_0_417), 
      .ZN(n_29));
   INV_X1 i_0_412 (.A(n_0_398), .ZN(n_0_397));
   OAI221_X1 i_0_413 (.A(n_0_399), .B1(n_0_408), .B2(n_0_407), .C1(n_0_502), 
      .C2(n_0_409), .ZN(n_0_398));
   AOI21_X1 i_0_414 (.A(n_0_400), .B1(n_0_479), .B2(n_0_406), .ZN(n_0_399));
   OAI21_X1 i_0_415 (.A(n_0_401), .B1(n_0_508), .B2(n_0_403), .ZN(n_0_400));
   NAND3_X1 i_0_416 (.A1(in_m[19]), .A2(n_0_484), .A3(n_0_402), .ZN(n_0_401));
   OAI21_X1 i_0_417 (.A(n_0_509), .B1(in_m[20]), .B2(n_0_505), .ZN(n_0_402));
   AOI21_X1 i_0_418 (.A(n_0_483), .B1(n_0_509), .B2(in_m[18]), .ZN(n_0_403));
   INV_X1 i_0_419 (.A(n_0_405), .ZN(n_0_404));
   NAND2_X1 i_0_420 (.A1(in_m[21]), .A2(n_0_484), .ZN(n_0_405));
   OAI33_X1 i_0_421 (.A1(in_m[19]), .A2(n_0_504), .A3(n_0_506), .B1(in_m[20]), 
      .B2(n_0_505), .B3(n_0_441), .ZN(n_0_406));
   NAND3_X1 i_0_422 (.A1(in_m[13]), .A2(n_0_474), .A3(n_0_477), .ZN(n_0_407));
   NAND2_X1 i_0_423 (.A1(n_0_504), .A2(in_m[15]), .ZN(n_0_408));
   AOI21_X1 i_0_424 (.A(n_0_412), .B1(in_m[12]), .B2(n_0_410), .ZN(n_0_409));
   INV_X1 i_0_425 (.A(n_0_411), .ZN(n_0_410));
   NAND2_X1 i_0_426 (.A1(n_0_503), .A2(n_0_471), .ZN(n_0_411));
   NOR3_X1 i_0_427 (.A1(n_0_504), .A2(n_0_478), .A3(n_0_476), .ZN(n_0_412));
   NAND3_X1 i_0_428 (.A1(n_0_502), .A2(in_m[11]), .A3(n_0_414), .ZN(n_0_413));
   OAI33_X1 i_0_429 (.A1(n_0_497), .A2(n_0_436), .A3(in_m[12]), .B1(in_m[16]), 
      .B2(n_0_472), .B3(n_0_501), .ZN(n_0_414));
   INV_X1 i_0_430 (.A(n_0_416), .ZN(n_0_415));
   NAND2_X1 i_0_431 (.A1(n_0_504), .A2(n_0_471), .ZN(n_0_416));
   AOI211_X1 i_0_432 (.A(n_0_420), .B(n_0_418), .C1(n_0_449), .C2(n_0_428), 
      .ZN(n_0_417));
   OAI21_X1 i_0_433 (.A(n_0_421), .B1(n_0_498), .B2(n_0_419), .ZN(n_0_418));
   AOI22_X1 i_0_434 (.A1(in_m[8]), .A2(n_0_426), .B1(n_0_501), .B2(in_m[12]), 
      .ZN(n_0_419));
   AOI211_X1 i_0_435 (.A(n_0_464), .B(n_0_452), .C1(n_0_496), .C2(n_0_430), 
      .ZN(n_0_420));
   NAND3_X1 i_0_436 (.A1(in_m[7]), .A2(n_0_422), .A3(n_0_424), .ZN(n_0_421));
   INV_X1 i_0_437 (.A(n_0_423), .ZN(n_0_422));
   NAND2_X1 i_0_438 (.A1(n_0_498), .A2(in_m[9]), .ZN(n_0_423));
   INV_X1 i_0_439 (.A(n_0_425), .ZN(n_0_424));
   NAND2_X1 i_0_440 (.A1(n_0_500), .A2(n_0_454), .ZN(n_0_425));
   INV_X1 i_0_441 (.A(n_0_427), .ZN(n_0_426));
   NAND2_X1 i_0_442 (.A1(n_0_499), .A2(n_0_454), .ZN(n_0_427));
   OR2_X1 i_0_443 (.A1(n_0_431), .A2(n_0_429), .ZN(n_0_428));
   OAI33_X1 i_0_444 (.A1(in_m[5]), .A2(n_0_490), .A3(n_0_430), .B1(in_m[10]), 
      .B2(n_0_495), .B3(n_0_493), .ZN(n_0_429));
   NAND3_X1 i_0_445 (.A1(n_0_495), .A2(in_m[4]), .A3(n_0_447), .ZN(n_0_430));
   AOI211_X1 i_0_446 (.A(n_0_491), .B(n_0_448), .C1(n_0_434), .C2(n_0_432), 
      .ZN(n_0_431));
   NAND3_X1 i_0_447 (.A1(in_m[1]), .A2(n_0_458), .A3(n_0_492), .ZN(n_0_432));
   INV_X1 i_0_448 (.A(n_0_434), .ZN(n_0_433));
   NAND2_X1 i_0_449 (.A1(n_0_494), .A2(in_m[5]), .ZN(n_0_434));
   INV_X1 i_0_450 (.A(n_0_436), .ZN(n_0_435));
   NAND2_X1 i_0_451 (.A1(n_0_473), .A2(n_0_438), .ZN(n_0_436));
   AND2_X1 i_0_452 (.A1(n_0_473), .A2(n_0_469), .ZN(n_0_437));
   AND2_X1 i_0_453 (.A1(n_0_477), .A2(n_0_469), .ZN(n_0_438));
   OAI21_X1 i_0_454 (.A(n_0_439), .B1(n_0_472), .B2(n_0_444), .ZN(n_30));
   AOI21_X1 i_0_455 (.A(n_0_440), .B1(n_0_482), .B2(n_0_443), .ZN(n_0_439));
   AOI221_X1 i_0_456 (.A(n_0_478), .B1(n_0_475), .B2(n_0_441), .C1(n_0_506), 
      .C2(n_0_442), .ZN(n_0_440));
   NAND2_X1 i_0_457 (.A1(n_0_506), .A2(in_m[15]), .ZN(n_0_441));
   NAND2_X1 i_0_458 (.A1(n_0_507), .A2(in_m[16]), .ZN(n_0_442));
   OAI21_X1 i_0_459 (.A(n_0_509), .B1(n_0_507), .B2(n_0_483), .ZN(n_0_443));
   AOI22_X1 i_0_460 (.A1(in_m[14]), .A2(n_0_470), .B1(n_0_469), .B2(n_0_445), 
      .ZN(n_0_444));
   OAI21_X1 i_0_461 (.A(n_0_446), .B1(n_0_465), .B2(n_0_462), .ZN(n_0_445));
   NAND3_X1 i_0_462 (.A1(n_0_449), .A2(n_0_447), .A3(n_0_456), .ZN(n_0_446));
   INV_X1 i_0_463 (.A(n_0_448), .ZN(n_0_447));
   NAND2_X1 i_0_464 (.A1(n_0_498), .A2(n_0_497), .ZN(n_0_448));
   INV_X1 i_0_465 (.A(n_0_450), .ZN(n_0_449));
   NAND2_X1 i_0_466 (.A1(n_0_496), .A2(n_0_451), .ZN(n_0_450));
   INV_X1 i_0_467 (.A(n_0_452), .ZN(n_0_451));
   NAND2_X1 i_0_468 (.A1(n_0_454), .A2(n_0_453), .ZN(n_0_452));
   NOR2_X1 i_0_469 (.A1(in_m[12]), .A2(in_m[11]), .ZN(n_0_453));
   INV_X1 i_0_470 (.A(n_0_455), .ZN(n_0_454));
   NAND2_X1 i_0_471 (.A1(n_0_502), .A2(n_0_501), .ZN(n_0_455));
   OAI21_X1 i_0_472 (.A(n_0_457), .B1(n_0_493), .B2(n_0_461), .ZN(n_0_456));
   NAND3_X1 i_0_473 (.A1(in_m[3]), .A2(n_0_458), .A3(n_0_460), .ZN(n_0_457));
   INV_X1 i_0_474 (.A(n_0_459), .ZN(n_0_458));
   NAND2_X1 i_0_475 (.A1(n_0_495), .A2(n_0_494), .ZN(n_0_459));
   OAI21_X1 i_0_476 (.A(n_0_492), .B1(in_m[5]), .B2(n_0_490), .ZN(n_0_460));
   AOI21_X1 i_0_477 (.A(in_m[6]), .B1(n_0_495), .B2(in_m[4]), .ZN(n_0_461));
   AOI211_X1 i_0_478 (.A(in_m[12]), .B(n_0_463), .C1(n_0_501), .C2(in_m[10]), 
      .ZN(n_0_462));
   AOI211_X1 i_0_479 (.A(in_m[13]), .B(in_m[11]), .C1(n_0_496), .C2(n_0_464), 
      .ZN(n_0_463));
   NAND2_X1 i_0_480 (.A1(n_0_497), .A2(in_m[6]), .ZN(n_0_464));
   AOI221_X1 i_0_481 (.A(in_m[13]), .B1(n_0_502), .B2(in_m[11]), .C1(n_0_468), 
      .C2(n_0_466), .ZN(n_0_465));
   INV_X1 i_0_482 (.A(n_0_467), .ZN(n_0_466));
   NAND2_X1 i_0_483 (.A1(n_0_502), .A2(n_0_500), .ZN(n_0_467));
   OAI21_X1 i_0_484 (.A(n_0_497), .B1(in_m[10]), .B2(n_0_495), .ZN(n_0_468));
   NOR2_X1 i_0_485 (.A1(in_m[16]), .A2(in_m[15]), .ZN(n_0_469));
   OAI21_X1 i_0_486 (.A(n_0_503), .B1(in_m[16]), .B2(n_0_501), .ZN(n_0_470));
   INV_X1 i_0_487 (.A(n_0_472), .ZN(n_0_471));
   NAND2_X1 i_0_488 (.A1(n_0_477), .A2(n_0_473), .ZN(n_0_472));
   NOR2_X1 i_0_489 (.A1(in_m[18]), .A2(n_0_476), .ZN(n_0_473));
   NOR2_X1 i_0_490 (.A1(in_m[19]), .A2(in_m[18]), .ZN(n_0_474));
   INV_X1 i_0_491 (.A(n_0_476), .ZN(n_0_475));
   NAND2_X1 i_0_492 (.A1(n_0_507), .A2(n_0_505), .ZN(n_0_476));
   INV_X1 i_0_493 (.A(n_0_478), .ZN(n_0_477));
   NAND2_X1 i_0_494 (.A1(n_0_509), .A2(n_0_481), .ZN(n_0_478));
   INV_X1 i_0_495 (.A(n_0_480), .ZN(n_0_479));
   NAND2_X1 i_0_496 (.A1(n_0_509), .A2(n_0_484), .ZN(n_0_480));
   INV_X1 i_0_497 (.A(n_0_482), .ZN(n_0_481));
   NAND2_X1 i_0_498 (.A1(n_0_508), .A2(n_0_484), .ZN(n_0_482));
   INV_X1 i_0_499 (.A(n_0_484), .ZN(n_0_483));
   NOR2_X1 i_0_500 (.A1(in_m[23]), .A2(in_m[22]), .ZN(n_0_484));
   INV_X1 i_0_501 (.A(n_0_14), .ZN(n_0_485));
   INV_X1 i_0_502 (.A(n_0_29), .ZN(n_0_486));
   INV_X1 i_0_503 (.A(n_0_12), .ZN(n_0_487));
   INV_X1 i_0_504 (.A(n_0_2), .ZN(n_0_488));
   INV_X1 i_0_505 (.A(in_m[1]), .ZN(n_0_489));
   INV_X1 i_0_506 (.A(in_m[2]), .ZN(n_0_490));
   INV_X1 i_0_507 (.A(in_m[3]), .ZN(n_0_491));
   INV_X1 i_0_508 (.A(in_m[4]), .ZN(n_0_492));
   INV_X1 i_0_509 (.A(in_m[5]), .ZN(n_0_493));
   INV_X1 i_0_510 (.A(in_m[6]), .ZN(n_0_494));
   INV_X1 i_0_511 (.A(in_m[7]), .ZN(n_0_495));
   INV_X1 i_0_512 (.A(in_m[8]), .ZN(n_0_496));
   INV_X1 i_0_513 (.A(in_m[9]), .ZN(n_0_497));
   INV_X1 i_0_514 (.A(in_m[10]), .ZN(n_0_498));
   INV_X1 i_0_515 (.A(in_m[11]), .ZN(n_0_499));
   INV_X1 i_0_516 (.A(in_m[12]), .ZN(n_0_500));
   INV_X1 i_0_517 (.A(in_m[13]), .ZN(n_0_501));
   INV_X1 i_0_518 (.A(in_m[14]), .ZN(n_0_502));
   INV_X1 i_0_519 (.A(in_m[15]), .ZN(n_0_503));
   INV_X1 i_0_520 (.A(in_m[16]), .ZN(n_0_504));
   INV_X1 i_0_521 (.A(in_m[17]), .ZN(n_0_505));
   INV_X1 i_0_522 (.A(in_m[18]), .ZN(n_0_506));
   INV_X1 i_0_523 (.A(in_m[19]), .ZN(n_0_507));
   INV_X1 i_0_524 (.A(in_m[20]), .ZN(n_0_508));
   INV_X1 i_0_525 (.A(in_m[21]), .ZN(n_0_509));
   INV_X1 i_0_526 (.A(in_e[0]), .ZN(n_0_510));
   INV_X1 i_0_527 (.A(in_e[1]), .ZN(n_0_511));
   INV_X1 i_0_528 (.A(in_e[2]), .ZN(n_0_512));
   INV_X1 i_0_529 (.A(in_e[3]), .ZN(n_0_513));
   INV_X1 i_0_530 (.A(in_e[6]), .ZN(n_0_514));
endmodule

module CLA_4bit__1_7(x, y, cO, s, p, g);
   input [3:0]x;
   input [3:0]y;
   input cO;
   output [3:0]s;
   output p;
   output g;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   FA_X1 i_0_0 (.A(1'b0), .B(x[0]), .CI(y[0]), .CO(n_0_0), .S(s[0]));
   FA_X1 i_0_1 (.A(y[1]), .B(x[1]), .CI(n_0_0), .CO(n_0_1), .S(s[1]));
   FA_X1 i_0_2 (.A(y[2]), .B(x[2]), .CI(n_0_1), .CO(n_0_2), .S(s[2]));
   AOI21_X1 i_0_3 (.A(n_0_5), .B1(n_0_3), .B2(n_0_4), .ZN(g));
   AOI22_X1 i_0_4 (.A1(y[3]), .A2(x[3]), .B1(x[2]), .B2(y[2]), .ZN(n_0_3));
   OAI211_X1 i_0_5 (.A(y[0]), .B(x[0]), .C1(x[2]), .C2(y[2]), .ZN(n_0_4));
   NOR2_X1 i_0_6 (.A1(y[3]), .A2(x[3]), .ZN(n_0_5));
   XNOR2_X1 i_0_7 (.A(y[3]), .B(n_0_6), .ZN(s[3]));
   XNOR2_X1 i_0_8 (.A(x[3]), .B(n_0_2), .ZN(n_0_6));
endmodule

module CLA_4bit__1_15(x, y, cO, s, p, g);
   input [3:0]x;
   input [3:0]y;
   input cO;
   output [3:0]s;
   output p;
   output g;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;

   FA_X1 i_0_0 (.A(cO), .B(x[0]), .CI(y[0]), .CO(n_0_0), .S(s[0]));
   FA_X1 i_0_1 (.A(y[1]), .B(x[1]), .CI(n_0_0), .CO(n_0_1), .S(s[1]));
   FA_X1 i_0_2 (.A(y[2]), .B(x[2]), .CI(n_0_1), .CO(n_0_2), .S(s[2]));
   OAI21_X1 i_0_3 (.A(n_0_4), .B1(n_0_3), .B2(n_0_6), .ZN(g));
   AOI22_X1 i_0_4 (.A1(y[2]), .A2(x[2]), .B1(x[0]), .B2(y[0]), .ZN(n_0_3));
   NAND2_X1 i_0_5 (.A1(y[3]), .A2(x[3]), .ZN(n_0_4));
   NOR2_X1 i_0_6 (.A1(n_0_6), .A2(n_0_5), .ZN(p));
   OAI22_X1 i_0_7 (.A1(y[1]), .A2(x[1]), .B1(x[0]), .B2(y[0]), .ZN(n_0_5));
   OAI22_X1 i_0_8 (.A1(y[3]), .A2(x[3]), .B1(x[2]), .B2(y[2]), .ZN(n_0_6));
   XNOR2_X1 i_0_9 (.A(y[3]), .B(n_0_7), .ZN(s[3]));
   XNOR2_X1 i_0_10 (.A(x[3]), .B(n_0_2), .ZN(n_0_7));
endmodule

module CLA_4bit__1_23(x, y, cO, s, p, g);
   input [3:0]x;
   input [3:0]y;
   input cO;
   output [3:0]s;
   output p;
   output g;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;

   FA_X1 i_0_0 (.A(cO), .B(x[0]), .CI(y[0]), .CO(n_0_0), .S(s[0]));
   FA_X1 i_0_1 (.A(y[1]), .B(x[1]), .CI(n_0_0), .CO(n_0_1), .S(s[1]));
   FA_X1 i_0_2 (.A(y[2]), .B(x[2]), .CI(n_0_1), .CO(n_0_2), .S(s[2]));
   OAI21_X1 i_0_3 (.A(n_0_4), .B1(n_0_3), .B2(n_0_6), .ZN(g));
   AOI22_X1 i_0_4 (.A1(y[2]), .A2(x[2]), .B1(x[0]), .B2(y[0]), .ZN(n_0_3));
   NAND2_X1 i_0_5 (.A1(y[3]), .A2(x[3]), .ZN(n_0_4));
   NOR2_X1 i_0_6 (.A1(n_0_6), .A2(n_0_5), .ZN(p));
   OAI22_X1 i_0_7 (.A1(y[1]), .A2(x[1]), .B1(x[0]), .B2(y[0]), .ZN(n_0_5));
   OAI22_X1 i_0_8 (.A1(y[3]), .A2(x[3]), .B1(x[2]), .B2(y[2]), .ZN(n_0_6));
   XNOR2_X1 i_0_9 (.A(y[3]), .B(n_0_7), .ZN(s[3]));
   XNOR2_X1 i_0_10 (.A(x[3]), .B(n_0_2), .ZN(n_0_7));
endmodule

module CLA_4bit__1_31(x, y, cO, s, p, g);
   input [3:0]x;
   input [3:0]y;
   input cO;
   output [3:0]s;
   output p;
   output g;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;

   FA_X1 i_0_0 (.A(cO), .B(x[0]), .CI(y[0]), .CO(n_0_0), .S(s[0]));
   FA_X1 i_0_1 (.A(y[1]), .B(x[1]), .CI(n_0_0), .CO(n_0_1), .S(s[1]));
   FA_X1 i_0_2 (.A(y[2]), .B(x[2]), .CI(n_0_1), .CO(n_0_2), .S(s[2]));
   OAI21_X1 i_0_3 (.A(n_0_4), .B1(n_0_3), .B2(n_0_6), .ZN(g));
   AOI22_X1 i_0_4 (.A1(y[2]), .A2(x[2]), .B1(x[0]), .B2(y[0]), .ZN(n_0_3));
   NAND2_X1 i_0_5 (.A1(y[3]), .A2(x[3]), .ZN(n_0_4));
   NOR2_X1 i_0_6 (.A1(n_0_6), .A2(n_0_5), .ZN(p));
   OAI22_X1 i_0_7 (.A1(y[1]), .A2(x[1]), .B1(x[0]), .B2(y[0]), .ZN(n_0_5));
   OAI22_X1 i_0_8 (.A1(y[3]), .A2(x[3]), .B1(x[2]), .B2(y[2]), .ZN(n_0_6));
   XNOR2_X1 i_0_9 (.A(y[3]), .B(n_0_7), .ZN(s[3]));
   XNOR2_X1 i_0_10 (.A(x[3]), .B(n_0_2), .ZN(n_0_7));
endmodule

module CLA_4bit__1_39(x, y, cO, s, p, g);
   input [3:0]x;
   input [3:0]y;
   input cO;
   output [3:0]s;
   output p;
   output g;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;

   FA_X1 i_0_0 (.A(cO), .B(x[0]), .CI(y[0]), .CO(n_0_0), .S(s[0]));
   FA_X1 i_0_1 (.A(y[1]), .B(x[1]), .CI(n_0_0), .CO(n_0_1), .S(s[1]));
   FA_X1 i_0_2 (.A(y[2]), .B(x[2]), .CI(n_0_1), .CO(n_0_2), .S(s[2]));
   OAI21_X1 i_0_3 (.A(n_0_4), .B1(n_0_3), .B2(n_0_6), .ZN(g));
   AOI22_X1 i_0_4 (.A1(y[2]), .A2(x[2]), .B1(x[0]), .B2(y[0]), .ZN(n_0_3));
   NAND2_X1 i_0_5 (.A1(y[3]), .A2(x[3]), .ZN(n_0_4));
   NOR2_X1 i_0_6 (.A1(n_0_6), .A2(n_0_5), .ZN(p));
   OAI22_X1 i_0_7 (.A1(y[1]), .A2(x[1]), .B1(x[0]), .B2(y[0]), .ZN(n_0_5));
   OAI22_X1 i_0_8 (.A1(y[3]), .A2(x[3]), .B1(x[2]), .B2(y[2]), .ZN(n_0_6));
   XNOR2_X1 i_0_9 (.A(y[3]), .B(n_0_7), .ZN(s[3]));
   XNOR2_X1 i_0_10 (.A(x[3]), .B(n_0_2), .ZN(n_0_7));
endmodule

module CLA_4bit(x, y, cO, s, p, g);
   input [3:0]x;
   input [3:0]y;
   input cO;
   output [3:0]s;
   output p;
   output g;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;

   FA_X1 i_0_0 (.A(cO), .B(x[0]), .CI(y[0]), .CO(n_0_0), .S(s[0]));
   FA_X1 i_0_1 (.A(y[1]), .B(x[1]), .CI(n_0_0), .CO(n_0_1), .S(s[1]));
   FA_X1 i_0_2 (.A(y[2]), .B(x[2]), .CI(n_0_1), .CO(n_0_2), .S(s[2]));
   OAI21_X1 i_0_3 (.A(n_0_4), .B1(n_0_3), .B2(n_0_6), .ZN(g));
   AOI22_X1 i_0_4 (.A1(y[2]), .A2(x[2]), .B1(x[0]), .B2(y[0]), .ZN(n_0_3));
   NAND2_X1 i_0_5 (.A1(y[3]), .A2(x[3]), .ZN(n_0_4));
   NOR2_X1 i_0_6 (.A1(n_0_6), .A2(n_0_5), .ZN(p));
   OAI22_X1 i_0_7 (.A1(y[1]), .A2(x[1]), .B1(x[0]), .B2(y[0]), .ZN(n_0_5));
   OAI22_X1 i_0_8 (.A1(y[3]), .A2(x[3]), .B1(x[2]), .B2(y[2]), .ZN(n_0_6));
   XNOR2_X1 i_0_9 (.A(y[3]), .B(n_0_7), .ZN(s[3]));
   XNOR2_X1 i_0_10 (.A(x[3]), .B(n_0_2), .ZN(n_0_7));
endmodule

module CLA_adder(A, B, Cin, Sum, Cout, Overflow);
   input [23:0]A;
   input [23:0]B;
   input Cin;
   output [23:0]Sum;
   output Cout;
   output Overflow;

   wire w_G;
   wire n_0_0;
   wire n_0_1;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   CLA_4bit__1_7 genblk1_0_stage1 (.x({A[3], A[2], A[1], A[0]}), .y({B[3], B[2], 
      B[1], B[0]}), .cO(), .s({Sum[3], Sum[2], Sum[1], Sum[0]}), .p(), .g(w_G));
   CLA_4bit__1_15 genblk1_1_stage1 (.x({A[7], A[6], A[5], A[4]}), .y({B[7], B[6], 
      B[5], B[4]}), .cO(w_G), .s({Sum[7], Sum[6], Sum[5], Sum[4]}), .p(n_1), 
      .g(n_0));
   CLA_4bit__1_23 genblk1_2_stage1 (.x({A[11], A[10], A[9], A[8]}), .y({B[11], 
      B[10], B[9], B[8]}), .cO(n_10), .s({Sum[11], Sum[10], Sum[9], Sum[8]}), 
      .p(n_3), .g(n_2));
   CLA_4bit__1_31 genblk1_3_stage1 (.x({A[15], A[14], A[13], A[12]}), .y({B[15], 
      B[14], B[13], B[12]}), .cO(n_11), .s({Sum[15], Sum[14], Sum[13], Sum[12]}), 
      .p(n_5), .g(n_4));
   CLA_4bit__1_39 genblk1_4_stage1 (.x({A[19], A[18], A[17], A[16]}), .y({B[19], 
      B[18], B[17], B[16]}), .cO(n_12), .s({Sum[19], Sum[18], Sum[17], Sum[16]}), 
      .p(n_7), .g(n_6));
   CLA_4bit genblk1_5_stage1 (.x({A[23], A[22], A[21], A[20]}), .y({B[23], B[22], 
      B[21], B[20]}), .cO(n_13), .s({Sum[23], Sum[22], Sum[21], Sum[20]}), 
      .p(n_9), .g(n_8));
   XOR2_X1 i_0_0 (.A(A[23]), .B(B[23]), .Z(n_0_0));
   XNOR2_X1 i_0_1 (.A(A[23]), .B(Sum[23]), .ZN(n_0_1));
   NOR2_X1 i_0_2 (.A1(n_0_0), .A2(n_0_1), .ZN(Overflow));
   AOI21_X1 i_1_0 (.A(n_0), .B1(n_1), .B2(w_G), .ZN(n_1_0));
   INV_X1 i_1_1 (.A(n_1_0), .ZN(n_10));
   AOI21_X1 i_1_2 (.A(n_2), .B1(n_3), .B2(n_10), .ZN(n_1_1));
   INV_X1 i_1_3 (.A(n_1_1), .ZN(n_11));
   AOI21_X1 i_1_4 (.A(n_4), .B1(n_5), .B2(n_11), .ZN(n_1_2));
   INV_X1 i_1_5 (.A(n_1_2), .ZN(n_12));
   AOI21_X1 i_1_6 (.A(n_6), .B1(n_7), .B2(n_12), .ZN(n_1_3));
   INV_X1 i_1_7 (.A(n_1_3), .ZN(n_13));
   AOI21_X1 i_1_8 (.A(n_8), .B1(n_9), .B2(n_13), .ZN(n_1_4));
   INV_X1 i_1_9 (.A(n_1_4), .ZN(Cout));
endmodule

module adder(a, b, out, of);
   input [31:0]a;
   input [31:0]b;
   output [31:0]out;
   output of;

   wire [24:0]o_m;
   wire [7:0]o_e;
   wire CLA_COUT;
   wire [23:0]CLA_SUM;
   wire [24:0]i_m;
   wire [7:0]i_e;
   wire n_0_6;
   wire n_0_0;
   wire n_0_7;
   wire n_0_1;
   wire n_0_8;
   wire n_0_2;
   wire n_0_9;
   wire n_0_3;
   wire n_0_10;
   wire n_0_4;
   wire n_0_11;
   wire n_0_5;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_317;
   wire n_0_318;
   wire n_0_319;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_332;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_337;
   wire n_0_338;
   wire n_0_339;
   wire n_0_340;
   wire n_0_341;
   wire n_0_342;
   wire n_0_343;
   wire n_0_344;
   wire n_0_345;
   wire n_0_346;
   wire n_0_347;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_355;
   wire n_0_356;
   wire n_0_357;
   wire n_0_358;
   wire n_0_359;
   wire n_0_360;
   wire n_0_361;
   wire n_0_362;
   wire n_0_363;
   wire n_0_364;
   wire n_0_365;
   wire n_0_366;
   wire n_0_367;
   wire n_0_368;
   wire n_0_369;
   wire n_0_370;
   wire n_0_371;
   wire n_0_372;
   wire n_0_373;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_377;
   wire n_0_378;
   wire n_0_379;
   wire n_0_380;
   wire n_0_381;
   wire n_0_382;
   wire n_0_383;
   wire n_0_384;
   wire n_0_385;
   wire n_0_386;
   wire n_0_387;
   wire n_0_388;
   wire n_0_389;
   wire n_0_390;
   wire n_0_391;
   wire n_0_392;
   wire n_0_393;
   wire n_0_394;
   wire n_0_395;
   wire n_0_396;
   wire n_0_397;
   wire n_0_398;
   wire n_0_399;
   wire n_0_400;
   wire n_0_401;
   wire n_0_402;
   wire n_0_403;
   wire n_0_404;
   wire n_0_405;
   wire n_0_406;
   wire n_0_407;
   wire n_0_408;
   wire n_0_409;
   wire n_0_410;
   wire n_0_411;
   wire n_0_412;
   wire n_0_413;
   wire n_0_414;
   wire n_0_415;
   wire n_0_416;
   wire n_0_417;
   wire n_0_418;
   wire n_0_419;
   wire n_0_420;
   wire n_0_421;
   wire n_0_422;
   wire n_0_423;
   wire n_0_424;
   wire n_0_425;
   wire n_0_426;
   wire n_0_427;
   wire n_0_428;
   wire n_0_429;
   wire n_0_430;
   wire n_0_431;
   wire n_0_432;
   wire n_0_433;
   wire n_0_434;
   wire n_0_435;
   wire n_0_436;
   wire n_0_437;
   wire n_0_438;
   wire n_0_439;
   wire n_0_440;
   wire n_0_441;
   wire n_0_442;
   wire n_0_443;
   wire n_0_444;
   wire n_0_445;
   wire n_0_446;
   wire n_0_447;
   wire n_0_448;
   wire n_0_449;
   wire n_0_450;
   wire n_0_451;
   wire n_0_452;
   wire n_0_453;
   wire n_0_454;
   wire n_0_455;
   wire n_0_456;
   wire n_0_457;
   wire n_0_458;
   wire n_0_459;
   wire n_0_460;
   wire n_0_461;
   wire n_0_462;
   wire n_0_463;
   wire n_0_464;
   wire n_0_465;
   wire n_0_466;
   wire n_0_467;
   wire n_0_468;
   wire n_0_469;
   wire n_0_470;
   wire n_0_471;
   wire n_0_472;
   wire n_0_473;
   wire n_0_474;
   wire n_0_475;
   wire n_0_476;
   wire n_0_477;
   wire n_0_478;
   wire n_0_479;
   wire n_0_480;
   wire n_0_481;
   wire n_0_482;
   wire n_0_483;
   wire n_0_484;
   wire n_0_485;
   wire n_0_486;
   wire n_0_487;
   wire n_0_488;
   wire n_0_489;
   wire n_0_490;
   wire n_0_491;
   wire n_0_492;
   wire n_0_493;
   wire n_0_494;
   wire n_0_495;
   wire n_0_496;
   wire n_0_497;
   wire n_0_498;
   wire n_0_499;
   wire n_0_500;
   wire n_0_501;
   wire n_0_502;
   wire n_0_503;
   wire n_0_504;
   wire n_0_505;
   wire n_0_506;
   wire n_0_507;
   wire n_0_508;
   wire n_0_509;
   wire n_0_510;
   wire n_0_511;
   wire n_0_512;
   wire n_0_513;
   wire n_0_514;
   wire n_0_515;
   wire n_0_516;
   wire n_0_517;
   wire n_0_518;
   wire n_0_519;
   wire n_0_520;
   wire n_0_521;
   wire n_0_522;
   wire n_0_523;
   wire n_0_524;
   wire n_0_525;
   wire n_0_526;
   wire n_0_527;
   wire n_0_528;
   wire n_0_529;
   wire n_0_530;
   wire n_0_531;
   wire n_0_532;
   wire n_0_533;
   wire n_0_534;
   wire n_0_535;
   wire n_0_536;

   addition_normaliser norm1 (.in_e(i_e), .in_m({uc_0, i_m[23], i_m[22], i_m[21], 
      i_m[20], i_m[19], i_m[18], i_m[17], i_m[16], i_m[15], i_m[14], i_m[13], 
      i_m[12], i_m[11], i_m[10], i_m[9], i_m[8], i_m[7], i_m[6], i_m[5], i_m[4], 
      i_m[3], i_m[2], i_m[1], i_m[0]}), .out_e(o_e), .out_m({uc_1, uc_2, o_m[22], 
      o_m[21], o_m[20], o_m[19], o_m[18], o_m[17], o_m[16], o_m[15], o_m[14], 
      o_m[13], o_m[12], o_m[11], o_m[10], o_m[9], o_m[8], o_m[7], o_m[6], o_m[5], 
      o_m[4], o_m[3], o_m[2], o_m[1], uc_3}));
   CLA_adder c1 (.A({n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, 
      n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0}), 
      .B({n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, 
      n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, n_24}), 
      .Cin(), .Sum(CLA_SUM), .Cout(CLA_COUT), .Overflow(of));
   DLH_X1 \i_m_reg[23]  (.D(CLA_SUM[23]), .G(n_48), .Q(i_m[23]));
   DLH_X1 \i_m_reg[22]  (.D(CLA_SUM[22]), .G(n_48), .Q(i_m[22]));
   DLH_X1 \i_m_reg[21]  (.D(CLA_SUM[21]), .G(n_48), .Q(i_m[21]));
   DLH_X1 \i_m_reg[20]  (.D(CLA_SUM[20]), .G(n_48), .Q(i_m[20]));
   DLH_X1 \i_m_reg[19]  (.D(CLA_SUM[19]), .G(n_48), .Q(i_m[19]));
   DLH_X1 \i_m_reg[18]  (.D(CLA_SUM[18]), .G(n_48), .Q(i_m[18]));
   DLH_X1 \i_m_reg[17]  (.D(CLA_SUM[17]), .G(n_48), .Q(i_m[17]));
   DLH_X1 \i_m_reg[16]  (.D(CLA_SUM[16]), .G(n_48), .Q(i_m[16]));
   DLH_X1 \i_m_reg[15]  (.D(CLA_SUM[15]), .G(n_48), .Q(i_m[15]));
   DLH_X1 \i_m_reg[14]  (.D(CLA_SUM[14]), .G(n_48), .Q(i_m[14]));
   DLH_X1 \i_m_reg[13]  (.D(CLA_SUM[13]), .G(n_48), .Q(i_m[13]));
   DLH_X1 \i_m_reg[12]  (.D(CLA_SUM[12]), .G(n_48), .Q(i_m[12]));
   DLH_X1 \i_m_reg[11]  (.D(CLA_SUM[11]), .G(n_48), .Q(i_m[11]));
   DLH_X1 \i_m_reg[10]  (.D(CLA_SUM[10]), .G(n_48), .Q(i_m[10]));
   DLH_X1 \i_m_reg[9]  (.D(CLA_SUM[9]), .G(n_48), .Q(i_m[9]));
   DLH_X1 \i_m_reg[8]  (.D(CLA_SUM[8]), .G(n_48), .Q(i_m[8]));
   DLH_X1 \i_m_reg[7]  (.D(CLA_SUM[7]), .G(n_48), .Q(i_m[7]));
   DLH_X1 \i_m_reg[6]  (.D(CLA_SUM[6]), .G(n_48), .Q(i_m[6]));
   DLH_X1 \i_m_reg[5]  (.D(CLA_SUM[5]), .G(n_48), .Q(i_m[5]));
   DLH_X1 \i_m_reg[4]  (.D(CLA_SUM[4]), .G(n_48), .Q(i_m[4]));
   DLH_X1 \i_m_reg[3]  (.D(CLA_SUM[3]), .G(n_48), .Q(i_m[3]));
   DLH_X1 \i_m_reg[2]  (.D(CLA_SUM[2]), .G(n_48), .Q(i_m[2]));
   DLH_X1 \i_m_reg[1]  (.D(CLA_SUM[1]), .G(n_48), .Q(i_m[1]));
   DLH_X1 \i_m_reg[0]  (.D(CLA_SUM[0]), .G(n_48), .Q(i_m[0]));
   DLH_X1 \i_e_reg[7]  (.D(n_56), .G(n_48), .Q(i_e[7]));
   DLH_X1 \i_e_reg[6]  (.D(n_55), .G(n_48), .Q(i_e[6]));
   DLH_X1 \i_e_reg[5]  (.D(n_54), .G(n_48), .Q(i_e[5]));
   DLH_X1 \i_e_reg[4]  (.D(n_53), .G(n_48), .Q(i_e[4]));
   DLH_X1 \i_e_reg[3]  (.D(n_52), .G(n_48), .Q(i_e[3]));
   DLH_X1 \i_e_reg[2]  (.D(n_51), .G(n_48), .Q(i_e[2]));
   DLH_X1 \i_e_reg[1]  (.D(n_50), .G(n_48), .Q(i_e[1]));
   DLH_X1 \i_e_reg[0]  (.D(n_49), .G(n_48), .Q(i_e[0]));
   HA_X1 i_0_0 (.A(n_50), .B(n_49), .CO(n_0_0), .S(n_0_6));
   HA_X1 i_0_1 (.A(n_51), .B(n_0_0), .CO(n_0_1), .S(n_0_7));
   HA_X1 i_0_2 (.A(n_52), .B(n_0_1), .CO(n_0_2), .S(n_0_8));
   HA_X1 i_0_3 (.A(n_53), .B(n_0_2), .CO(n_0_3), .S(n_0_9));
   HA_X1 i_0_4 (.A(n_54), .B(n_0_3), .CO(n_0_4), .S(n_0_10));
   HA_X1 i_0_5 (.A(n_55), .B(n_0_4), .CO(n_0_5), .S(n_0_11));
   OAI21_X1 i_0_6 (.A(n_0_12), .B1(a[0]), .B2(n_0_397), .ZN(n_0));
   AOI22_X1 i_0_7 (.A1(a[0]), .A2(n_0_394), .B1(b[0]), .B2(n_0_437), .ZN(n_0_12));
   OAI21_X1 i_0_8 (.A(n_0_13), .B1(a[1]), .B2(n_0_397), .ZN(n_1));
   AOI22_X1 i_0_9 (.A1(a[1]), .A2(n_0_394), .B1(b[1]), .B2(n_0_437), .ZN(n_0_13));
   OAI222_X1 i_0_10 (.A1(n_0_509), .A2(n_0_438), .B1(a[2]), .B2(n_0_397), 
      .C1(n_0_480), .C2(n_0_395), .ZN(n_2));
   OAI21_X1 i_0_11 (.A(n_0_14), .B1(a[3]), .B2(n_0_397), .ZN(n_3));
   AOI22_X1 i_0_12 (.A1(a[3]), .A2(n_0_394), .B1(b[3]), .B2(n_0_437), .ZN(n_0_14));
   OAI222_X1 i_0_13 (.A1(n_0_511), .A2(n_0_438), .B1(a[4]), .B2(n_0_397), 
      .C1(n_0_481), .C2(n_0_395), .ZN(n_4));
   OAI21_X1 i_0_14 (.A(n_0_15), .B1(a[5]), .B2(n_0_397), .ZN(n_5));
   AOI22_X1 i_0_15 (.A1(a[5]), .A2(n_0_394), .B1(b[5]), .B2(n_0_437), .ZN(n_0_15));
   OAI222_X1 i_0_16 (.A1(n_0_513), .A2(n_0_438), .B1(a[6]), .B2(n_0_397), 
      .C1(n_0_482), .C2(n_0_395), .ZN(n_6));
   OAI222_X1 i_0_17 (.A1(n_0_514), .A2(n_0_438), .B1(a[7]), .B2(n_0_397), 
      .C1(n_0_483), .C2(n_0_395), .ZN(n_7));
   OAI222_X1 i_0_18 (.A1(n_0_515), .A2(n_0_438), .B1(a[8]), .B2(n_0_397), 
      .C1(n_0_484), .C2(n_0_395), .ZN(n_8));
   OAI222_X1 i_0_19 (.A1(n_0_516), .A2(n_0_438), .B1(a[9]), .B2(n_0_397), 
      .C1(n_0_485), .C2(n_0_395), .ZN(n_9));
   OAI222_X1 i_0_20 (.A1(n_0_517), .A2(n_0_438), .B1(a[10]), .B2(n_0_397), 
      .C1(n_0_486), .C2(n_0_395), .ZN(n_10));
   OAI222_X1 i_0_21 (.A1(n_0_518), .A2(n_0_438), .B1(a[11]), .B2(n_0_397), 
      .C1(n_0_487), .C2(n_0_395), .ZN(n_11));
   OAI222_X1 i_0_22 (.A1(n_0_519), .A2(n_0_438), .B1(a[12]), .B2(n_0_397), 
      .C1(n_0_488), .C2(n_0_395), .ZN(n_12));
   OAI222_X1 i_0_23 (.A1(n_0_520), .A2(n_0_438), .B1(a[13]), .B2(n_0_397), 
      .C1(n_0_489), .C2(n_0_395), .ZN(n_13));
   OAI222_X1 i_0_24 (.A1(n_0_521), .A2(n_0_438), .B1(a[14]), .B2(n_0_397), 
      .C1(n_0_490), .C2(n_0_395), .ZN(n_14));
   OAI222_X1 i_0_25 (.A1(n_0_522), .A2(n_0_438), .B1(a[15]), .B2(n_0_397), 
      .C1(n_0_491), .C2(n_0_395), .ZN(n_15));
   OAI21_X1 i_0_26 (.A(n_0_16), .B1(n_0_492), .B2(n_0_395), .ZN(n_16));
   AOI22_X1 i_0_27 (.A1(b[16]), .A2(n_0_437), .B1(n_0_492), .B2(n_0_396), 
      .ZN(n_0_16));
   OAI222_X1 i_0_28 (.A1(n_0_523), .A2(n_0_438), .B1(a[17]), .B2(n_0_397), 
      .C1(n_0_493), .C2(n_0_395), .ZN(n_17));
   OAI222_X1 i_0_29 (.A1(n_0_524), .A2(n_0_438), .B1(a[18]), .B2(n_0_397), 
      .C1(n_0_494), .C2(n_0_395), .ZN(n_18));
   OAI222_X1 i_0_30 (.A1(n_0_525), .A2(n_0_438), .B1(a[19]), .B2(n_0_397), 
      .C1(n_0_495), .C2(n_0_395), .ZN(n_19));
   OAI222_X1 i_0_31 (.A1(n_0_526), .A2(n_0_438), .B1(a[20]), .B2(n_0_397), 
      .C1(n_0_496), .C2(n_0_395), .ZN(n_20));
   OAI222_X1 i_0_32 (.A1(n_0_527), .A2(n_0_438), .B1(a[21]), .B2(n_0_397), 
      .C1(n_0_497), .C2(n_0_395), .ZN(n_21));
   OAI222_X1 i_0_33 (.A1(n_0_528), .A2(n_0_438), .B1(a[22]), .B2(n_0_397), 
      .C1(n_0_498), .C2(n_0_395), .ZN(n_22));
   OAI221_X1 i_0_34 (.A(n_0_438), .B1(n_0_404), .B2(n_0_397), .C1(n_0_405), 
      .C2(n_0_396), .ZN(n_23));
   OAI21_X1 i_0_35 (.A(n_0_17), .B1(b[0]), .B2(n_0_356), .ZN(n_24));
   AOI21_X1 i_0_36 (.A(n_0_18), .B1(b[0]), .B2(n_0_350), .ZN(n_0_17));
   OAI221_X1 i_0_37 (.A(n_0_19), .B1(n_0_301), .B2(n_0_24), .C1(n_0_306), 
      .C2(n_0_20), .ZN(n_0_18));
   AOI22_X1 i_0_38 (.A1(n_0_352), .A2(n_0_24), .B1(n_0_353), .B2(n_0_20), 
      .ZN(n_0_19));
   AOI22_X1 i_0_39 (.A1(n_0_254), .A2(n_0_32), .B1(n_0_22), .B2(n_0_21), 
      .ZN(n_0_20));
   AOI21_X1 i_0_40 (.A(n_0_272), .B1(n_0_309), .B2(n_0_52), .ZN(n_0_21));
   OAI221_X1 i_0_41 (.A(n_0_310), .B1(n_0_323), .B2(n_0_23), .C1(n_0_322), 
      .C2(n_0_81), .ZN(n_0_22));
   AOI222_X1 i_0_42 (.A1(a[16]), .A2(n_0_117), .B1(a[0]), .B2(n_0_317), .C1(a[8]), 
      .C2(n_0_232), .ZN(n_0_23));
   AOI22_X1 i_0_43 (.A1(n_0_261), .A2(n_0_37), .B1(n_0_26), .B2(n_0_25), 
      .ZN(n_0_24));
   AOI21_X1 i_0_44 (.A(n_0_281), .B1(n_0_326), .B2(n_0_47), .ZN(n_0_25));
   OAI221_X1 i_0_45 (.A(n_0_327), .B1(n_0_335), .B2(n_0_27), .C1(n_0_334), 
      .C2(n_0_75), .ZN(n_0_26));
   AOI222_X1 i_0_46 (.A1(b[8]), .A2(n_0_226), .B1(b[16]), .B2(n_0_124), .C1(b[0]), 
      .C2(n_0_330), .ZN(n_0_27));
   OAI211_X1 i_0_47 (.A(n_0_29), .B(n_0_28), .C1(b[1]), .C2(n_0_356), .ZN(n_25));
   AOI22_X1 i_0_48 (.A1(b[1]), .A2(n_0_350), .B1(n_0_353), .B2(n_0_31), .ZN(
      n_0_28));
   AOI21_X1 i_0_49 (.A(n_0_30), .B1(n_0_352), .B2(n_0_36), .ZN(n_0_29));
   OAI22_X1 i_0_50 (.A1(n_0_301), .A2(n_0_36), .B1(n_0_306), .B2(n_0_31), 
      .ZN(n_0_30));
   AOI22_X1 i_0_51 (.A1(n_0_271), .A2(n_0_32), .B1(n_0_254), .B2(n_0_51), 
      .ZN(n_0_31));
   INV_X1 i_0_52 (.A(n_0_33), .ZN(n_0_32));
   AOI21_X1 i_0_53 (.A(n_0_34), .B1(n_0_309), .B2(n_0_61), .ZN(n_0_33));
   AOI221_X1 i_0_54 (.A(n_0_309), .B1(n_0_322), .B2(n_0_35), .C1(n_0_323), 
      .C2(n_0_95), .ZN(n_0_34));
   AOI222_X1 i_0_55 (.A1(a[1]), .A2(n_0_317), .B1(a[17]), .B2(n_0_117), .C1(a[9]), 
      .C2(n_0_232), .ZN(n_0_35));
   AOI22_X1 i_0_56 (.A1(n_0_261), .A2(n_0_45), .B1(n_0_280), .B2(n_0_37), 
      .ZN(n_0_36));
   AOI21_X1 i_0_57 (.A(n_0_38), .B1(n_0_326), .B2(n_0_65), .ZN(n_0_37));
   AOI221_X1 i_0_58 (.A(n_0_326), .B1(n_0_334), .B2(n_0_39), .C1(n_0_335), 
      .C2(n_0_89), .ZN(n_0_38));
   INV_X1 i_0_59 (.A(n_0_40), .ZN(n_0_39));
   AOI222_X1 i_0_60 (.A1(b[1]), .A2(n_0_330), .B1(b[17]), .B2(n_0_124), .C1(b[9]), 
      .C2(n_0_226), .ZN(n_0_40));
   OAI21_X1 i_0_61 (.A(n_0_41), .B1(b[2]), .B2(n_0_356), .ZN(n_26));
   AOI21_X1 i_0_62 (.A(n_0_42), .B1(b[2]), .B2(n_0_350), .ZN(n_0_41));
   OAI221_X1 i_0_63 (.A(n_0_43), .B1(n_0_306), .B2(n_0_50), .C1(n_0_301), 
      .C2(n_0_44), .ZN(n_0_42));
   AOI22_X1 i_0_64 (.A1(n_0_352), .A2(n_0_44), .B1(n_0_353), .B2(n_0_50), 
      .ZN(n_0_43));
   AOI22_X1 i_0_65 (.A1(n_0_280), .A2(n_0_45), .B1(n_0_261), .B2(n_0_64), 
      .ZN(n_0_44));
   OAI21_X1 i_0_66 (.A(n_0_46), .B1(n_0_326), .B2(n_0_47), .ZN(n_0_45));
   NAND2_X1 i_0_67 (.A1(n_0_326), .A2(n_0_74), .ZN(n_0_46));
   INV_X1 i_0_68 (.A(n_0_48), .ZN(n_0_47));
   AOI22_X1 i_0_69 (.A1(n_0_334), .A2(n_0_49), .B1(n_0_335), .B2(n_0_103), 
      .ZN(n_0_48));
   AOI222_X1 i_0_70 (.A1(b[18]), .A2(n_0_124), .B1(b[2]), .B2(n_0_330), .C1(
      b[10]), .C2(n_0_226), .ZN(n_0_49));
   AOI22_X1 i_0_71 (.A1(n_0_254), .A2(n_0_59), .B1(n_0_271), .B2(n_0_51), 
      .ZN(n_0_50));
   AOI22_X1 i_0_72 (.A1(n_0_310), .A2(n_0_52), .B1(n_0_309), .B2(n_0_79), 
      .ZN(n_0_51));
   INV_X1 i_0_73 (.A(n_0_53), .ZN(n_0_52));
   AOI22_X1 i_0_74 (.A1(n_0_323), .A2(n_0_108), .B1(n_0_322), .B2(n_0_54), 
      .ZN(n_0_53));
   AOI222_X1 i_0_75 (.A1(a[10]), .A2(n_0_232), .B1(a[18]), .B2(n_0_117), 
      .C1(a[2]), .C2(n_0_317), .ZN(n_0_54));
   OAI21_X1 i_0_76 (.A(n_0_55), .B1(b[3]), .B2(n_0_356), .ZN(n_27));
   AOI21_X1 i_0_77 (.A(n_0_56), .B1(b[3]), .B2(n_0_350), .ZN(n_0_55));
   OAI221_X1 i_0_78 (.A(n_0_57), .B1(n_0_301), .B2(n_0_63), .C1(n_0_306), 
      .C2(n_0_58), .ZN(n_0_56));
   AOI22_X1 i_0_79 (.A1(n_0_352), .A2(n_0_63), .B1(n_0_353), .B2(n_0_58), 
      .ZN(n_0_57));
   AOI22_X1 i_0_80 (.A1(n_0_254), .A2(n_0_78), .B1(n_0_271), .B2(n_0_59), 
      .ZN(n_0_58));
   AOI21_X1 i_0_81 (.A(n_0_60), .B1(n_0_309), .B2(n_0_93), .ZN(n_0_59));
   NOR2_X1 i_0_82 (.A1(n_0_309), .A2(n_0_61), .ZN(n_0_60));
   AOI22_X1 i_0_83 (.A1(n_0_323), .A2(n_0_116), .B1(n_0_322), .B2(n_0_62), 
      .ZN(n_0_61));
   AOI222_X1 i_0_84 (.A1(a[11]), .A2(n_0_232), .B1(a[19]), .B2(n_0_117), 
      .C1(a[3]), .C2(n_0_317), .ZN(n_0_62));
   AOI22_X1 i_0_85 (.A1(n_0_261), .A2(n_0_72), .B1(n_0_280), .B2(n_0_64), 
      .ZN(n_0_63));
   AOI22_X1 i_0_86 (.A1(n_0_327), .A2(n_0_65), .B1(n_0_326), .B2(n_0_87), 
      .ZN(n_0_64));
   INV_X1 i_0_87 (.A(n_0_66), .ZN(n_0_65));
   AOI22_X1 i_0_88 (.A1(n_0_335), .A2(n_0_123), .B1(n_0_334), .B2(n_0_67), 
      .ZN(n_0_66));
   AOI222_X1 i_0_89 (.A1(b[11]), .A2(n_0_226), .B1(b[3]), .B2(n_0_330), .C1(
      b[19]), .C2(n_0_124), .ZN(n_0_67));
   OAI21_X1 i_0_90 (.A(n_0_68), .B1(n_0_354), .B2(n_0_76), .ZN(n_28));
   AOI21_X1 i_0_91 (.A(n_0_69), .B1(n_0_305), .B2(n_0_76), .ZN(n_0_68));
   OAI221_X1 i_0_92 (.A(n_0_70), .B1(n_0_301), .B2(n_0_71), .C1(b[4]), .C2(
      n_0_356), .ZN(n_0_69));
   AOI22_X1 i_0_93 (.A1(b[4]), .A2(n_0_350), .B1(n_0_352), .B2(n_0_71), .ZN(
      n_0_70));
   AOI22_X1 i_0_94 (.A1(n_0_261), .A2(n_0_86), .B1(n_0_280), .B2(n_0_72), 
      .ZN(n_0_71));
   AOI21_X1 i_0_95 (.A(n_0_73), .B1(n_0_326), .B2(n_0_101), .ZN(n_0_72));
   NOR2_X1 i_0_96 (.A1(n_0_326), .A2(n_0_74), .ZN(n_0_73));
   AOI22_X1 i_0_97 (.A1(n_0_334), .A2(n_0_75), .B1(n_0_335), .B2(n_0_137), 
      .ZN(n_0_74));
   AOI222_X1 i_0_98 (.A1(b[12]), .A2(n_0_226), .B1(b[20]), .B2(n_0_124), 
      .C1(b[4]), .C2(n_0_330), .ZN(n_0_75));
   INV_X1 i_0_99 (.A(n_0_77), .ZN(n_0_76));
   AOI22_X1 i_0_100 (.A1(n_0_254), .A2(n_0_92), .B1(n_0_271), .B2(n_0_78), 
      .ZN(n_0_77));
   AOI22_X1 i_0_101 (.A1(n_0_310), .A2(n_0_79), .B1(n_0_309), .B2(n_0_106), 
      .ZN(n_0_78));
   INV_X1 i_0_102 (.A(n_0_80), .ZN(n_0_79));
   AOI22_X1 i_0_103 (.A1(n_0_323), .A2(n_0_132), .B1(n_0_322), .B2(n_0_81), 
      .ZN(n_0_80));
   AOI222_X1 i_0_104 (.A1(a[12]), .A2(n_0_232), .B1(a[20]), .B2(n_0_117), 
      .C1(a[4]), .C2(n_0_317), .ZN(n_0_81));
   OAI21_X1 i_0_105 (.A(n_0_82), .B1(b[5]), .B2(n_0_356), .ZN(n_29));
   AOI21_X1 i_0_106 (.A(n_0_83), .B1(b[5]), .B2(n_0_350), .ZN(n_0_82));
   OAI221_X1 i_0_107 (.A(n_0_84), .B1(n_0_306), .B2(n_0_91), .C1(n_0_301), 
      .C2(n_0_85), .ZN(n_0_83));
   AOI22_X1 i_0_108 (.A1(n_0_353), .A2(n_0_91), .B1(n_0_352), .B2(n_0_85), 
      .ZN(n_0_84));
   AOI22_X1 i_0_109 (.A1(n_0_261), .A2(n_0_100), .B1(n_0_280), .B2(n_0_86), 
      .ZN(n_0_85));
   AOI22_X1 i_0_110 (.A1(n_0_327), .A2(n_0_87), .B1(n_0_326), .B2(n_0_121), 
      .ZN(n_0_86));
   OAI21_X1 i_0_111 (.A(n_0_88), .B1(n_0_335), .B2(n_0_89), .ZN(n_0_87));
   NAND2_X1 i_0_112 (.A1(n_0_335), .A2(n_0_150), .ZN(n_0_88));
   INV_X1 i_0_113 (.A(n_0_90), .ZN(n_0_89));
   AOI222_X1 i_0_114 (.A1(b[13]), .A2(n_0_226), .B1(b[21]), .B2(n_0_124), 
      .C1(b[5]), .C2(n_0_330), .ZN(n_0_90));
   AOI22_X1 i_0_115 (.A1(n_0_254), .A2(n_0_105), .B1(n_0_271), .B2(n_0_92), 
      .ZN(n_0_91));
   AOI22_X1 i_0_116 (.A1(n_0_310), .A2(n_0_93), .B1(n_0_309), .B2(n_0_114), 
      .ZN(n_0_92));
   INV_X1 i_0_117 (.A(n_0_94), .ZN(n_0_93));
   AOI22_X1 i_0_118 (.A1(n_0_322), .A2(n_0_95), .B1(n_0_323), .B2(n_0_145), 
      .ZN(n_0_94));
   AOI222_X1 i_0_119 (.A1(a[13]), .A2(n_0_232), .B1(a[21]), .B2(n_0_117), 
      .C1(a[5]), .C2(n_0_317), .ZN(n_0_95));
   OAI21_X1 i_0_120 (.A(n_0_96), .B1(b[6]), .B2(n_0_356), .ZN(n_30));
   AOI21_X1 i_0_121 (.A(n_0_97), .B1(b[6]), .B2(n_0_350), .ZN(n_0_96));
   OAI221_X1 i_0_122 (.A(n_0_98), .B1(n_0_301), .B2(n_0_99), .C1(n_0_306), 
      .C2(n_0_104), .ZN(n_0_97));
   AOI22_X1 i_0_123 (.A1(n_0_353), .A2(n_0_104), .B1(n_0_352), .B2(n_0_99), 
      .ZN(n_0_98));
   AOI22_X1 i_0_124 (.A1(n_0_261), .A2(n_0_119), .B1(n_0_280), .B2(n_0_100), 
      .ZN(n_0_99));
   AOI22_X1 i_0_125 (.A1(n_0_326), .A2(n_0_135), .B1(n_0_327), .B2(n_0_101), 
      .ZN(n_0_100));
   INV_X1 i_0_126 (.A(n_0_102), .ZN(n_0_101));
   AOI22_X1 i_0_127 (.A1(n_0_334), .A2(n_0_103), .B1(n_0_335), .B2(n_0_164), 
      .ZN(n_0_102));
   AOI222_X1 i_0_128 (.A1(b[14]), .A2(n_0_226), .B1(b[22]), .B2(n_0_124), 
      .C1(b[6]), .C2(n_0_330), .ZN(n_0_103));
   AOI22_X1 i_0_129 (.A1(n_0_254), .A2(n_0_113), .B1(n_0_271), .B2(n_0_105), 
      .ZN(n_0_104));
   AOI22_X1 i_0_130 (.A1(n_0_310), .A2(n_0_106), .B1(n_0_309), .B2(n_0_130), 
      .ZN(n_0_105));
   INV_X1 i_0_131 (.A(n_0_107), .ZN(n_0_106));
   AOI22_X1 i_0_132 (.A1(n_0_323), .A2(n_0_159), .B1(n_0_322), .B2(n_0_108), 
      .ZN(n_0_107));
   AOI222_X1 i_0_133 (.A1(a[14]), .A2(n_0_232), .B1(a[22]), .B2(n_0_117), 
      .C1(a[6]), .C2(n_0_317), .ZN(n_0_108));
   OAI21_X1 i_0_134 (.A(n_0_109), .B1(b[7]), .B2(n_0_356), .ZN(n_31));
   AOI21_X1 i_0_135 (.A(n_0_110), .B1(b[7]), .B2(n_0_350), .ZN(n_0_109));
   OAI221_X1 i_0_136 (.A(n_0_111), .B1(n_0_306), .B2(n_0_112), .C1(n_0_301), 
      .C2(n_0_118), .ZN(n_0_110));
   AOI22_X1 i_0_137 (.A1(n_0_352), .A2(n_0_118), .B1(n_0_353), .B2(n_0_112), 
      .ZN(n_0_111));
   AOI22_X1 i_0_138 (.A1(n_0_271), .A2(n_0_113), .B1(n_0_254), .B2(n_0_129), 
      .ZN(n_0_112));
   AOI22_X1 i_0_139 (.A1(n_0_310), .A2(n_0_114), .B1(n_0_309), .B2(n_0_143), 
      .ZN(n_0_113));
   INV_X1 i_0_140 (.A(n_0_115), .ZN(n_0_114));
   AOI22_X1 i_0_141 (.A1(n_0_323), .A2(n_0_178), .B1(n_0_322), .B2(n_0_116), 
      .ZN(n_0_115));
   AOI222_X1 i_0_142 (.A1(n_0_404), .A2(n_0_117), .B1(a[7]), .B2(n_0_317), 
      .C1(a[15]), .C2(n_0_232), .ZN(n_0_116));
   NOR2_X1 i_0_143 (.A1(n_0_321), .A2(n_0_319), .ZN(n_0_117));
   AOI22_X1 i_0_144 (.A1(n_0_280), .A2(n_0_119), .B1(n_0_261), .B2(n_0_134), 
      .ZN(n_0_118));
   OAI21_X1 i_0_145 (.A(n_0_120), .B1(n_0_326), .B2(n_0_121), .ZN(n_0_119));
   NAND2_X1 i_0_146 (.A1(n_0_326), .A2(n_0_149), .ZN(n_0_120));
   INV_X1 i_0_147 (.A(n_0_122), .ZN(n_0_121));
   OAI22_X1 i_0_148 (.A1(n_0_334), .A2(n_0_173), .B1(n_0_335), .B2(n_0_123), 
      .ZN(n_0_122));
   AOI222_X1 i_0_149 (.A1(b[15]), .A2(n_0_226), .B1(b[7]), .B2(n_0_330), 
      .C1(n_0_402), .C2(n_0_124), .ZN(n_0_123));
   NOR2_X1 i_0_150 (.A1(n_0_333), .A2(n_0_332), .ZN(n_0_124));
   OAI21_X1 i_0_151 (.A(n_0_125), .B1(b[8]), .B2(n_0_356), .ZN(n_32));
   AOI21_X1 i_0_152 (.A(n_0_126), .B1(b[8]), .B2(n_0_350), .ZN(n_0_125));
   OAI221_X1 i_0_153 (.A(n_0_127), .B1(n_0_306), .B2(n_0_128), .C1(n_0_301), 
      .C2(n_0_133), .ZN(n_0_126));
   AOI22_X1 i_0_154 (.A1(n_0_352), .A2(n_0_133), .B1(n_0_353), .B2(n_0_128), 
      .ZN(n_0_127));
   AOI22_X1 i_0_155 (.A1(n_0_254), .A2(n_0_142), .B1(n_0_271), .B2(n_0_129), 
      .ZN(n_0_128));
   AOI22_X1 i_0_156 (.A1(n_0_310), .A2(n_0_130), .B1(n_0_309), .B2(n_0_157), 
      .ZN(n_0_129));
   INV_X1 i_0_157 (.A(n_0_131), .ZN(n_0_130));
   AOI22_X1 i_0_158 (.A1(n_0_322), .A2(n_0_132), .B1(n_0_323), .B2(n_0_186), 
      .ZN(n_0_131));
   AOI22_X1 i_0_159 (.A1(a[8]), .A2(n_0_317), .B1(a[16]), .B2(n_0_232), .ZN(
      n_0_132));
   AOI22_X1 i_0_160 (.A1(n_0_261), .A2(n_0_147), .B1(n_0_280), .B2(n_0_134), 
      .ZN(n_0_133));
   AOI22_X1 i_0_161 (.A1(n_0_327), .A2(n_0_135), .B1(n_0_326), .B2(n_0_162), 
      .ZN(n_0_134));
   OAI21_X1 i_0_162 (.A(n_0_136), .B1(n_0_334), .B2(n_0_191), .ZN(n_0_135));
   NAND2_X1 i_0_163 (.A1(n_0_334), .A2(n_0_137), .ZN(n_0_136));
   AOI22_X1 i_0_164 (.A1(b[8]), .A2(n_0_330), .B1(b[16]), .B2(n_0_226), .ZN(
      n_0_137));
   OAI211_X1 i_0_165 (.A(n_0_138), .B(n_0_140), .C1(b[9]), .C2(n_0_356), 
      .ZN(n_33));
   AOI21_X1 i_0_166 (.A(n_0_139), .B1(n_0_353), .B2(n_0_141), .ZN(n_0_138));
   OAI22_X1 i_0_167 (.A1(n_0_301), .A2(n_0_146), .B1(n_0_306), .B2(n_0_141), 
      .ZN(n_0_139));
   AOI22_X1 i_0_168 (.A1(b[9]), .A2(n_0_350), .B1(n_0_352), .B2(n_0_146), 
      .ZN(n_0_140));
   AOI22_X1 i_0_169 (.A1(n_0_271), .A2(n_0_142), .B1(n_0_254), .B2(n_0_155), 
      .ZN(n_0_141));
   AOI22_X1 i_0_170 (.A1(n_0_310), .A2(n_0_143), .B1(n_0_309), .B2(n_0_176), 
      .ZN(n_0_142));
   OAI21_X1 i_0_171 (.A(n_0_144), .B1(n_0_322), .B2(n_0_199), .ZN(n_0_143));
   NAND2_X1 i_0_172 (.A1(n_0_322), .A2(n_0_145), .ZN(n_0_144));
   AOI22_X1 i_0_173 (.A1(a[9]), .A2(n_0_317), .B1(a[17]), .B2(n_0_232), .ZN(
      n_0_145));
   AOI22_X1 i_0_174 (.A1(n_0_261), .A2(n_0_161), .B1(n_0_280), .B2(n_0_147), 
      .ZN(n_0_146));
   AOI21_X1 i_0_175 (.A(n_0_148), .B1(n_0_326), .B2(n_0_171), .ZN(n_0_147));
   NOR2_X1 i_0_176 (.A1(n_0_326), .A2(n_0_149), .ZN(n_0_148));
   AOI22_X1 i_0_177 (.A1(n_0_334), .A2(n_0_150), .B1(n_0_335), .B2(n_0_204), 
      .ZN(n_0_149));
   AOI22_X1 i_0_178 (.A1(b[9]), .A2(n_0_330), .B1(b[17]), .B2(n_0_226), .ZN(
      n_0_150));
   OAI21_X1 i_0_179 (.A(n_0_151), .B1(b[10]), .B2(n_0_356), .ZN(n_34));
   AOI21_X1 i_0_180 (.A(n_0_152), .B1(b[10]), .B2(n_0_350), .ZN(n_0_151));
   OAI221_X1 i_0_181 (.A(n_0_153), .B1(n_0_301), .B2(n_0_160), .C1(n_0_306), 
      .C2(n_0_154), .ZN(n_0_152));
   AOI22_X1 i_0_182 (.A1(n_0_352), .A2(n_0_160), .B1(n_0_353), .B2(n_0_154), 
      .ZN(n_0_153));
   AOI22_X1 i_0_183 (.A1(n_0_254), .A2(n_0_175), .B1(n_0_271), .B2(n_0_155), 
      .ZN(n_0_154));
   OAI21_X1 i_0_184 (.A(n_0_156), .B1(n_0_309), .B2(n_0_157), .ZN(n_0_155));
   NAND2_X1 i_0_185 (.A1(n_0_309), .A2(n_0_185), .ZN(n_0_156));
   AOI21_X1 i_0_186 (.A(n_0_158), .B1(n_0_323), .B2(n_0_217), .ZN(n_0_157));
   NOR2_X1 i_0_187 (.A1(n_0_323), .A2(n_0_159), .ZN(n_0_158));
   AOI22_X1 i_0_188 (.A1(a[10]), .A2(n_0_317), .B1(a[18]), .B2(n_0_232), 
      .ZN(n_0_159));
   AOI22_X1 i_0_189 (.A1(n_0_261), .A2(n_0_169), .B1(n_0_280), .B2(n_0_161), 
      .ZN(n_0_160));
   AOI22_X1 i_0_190 (.A1(n_0_326), .A2(n_0_190), .B1(n_0_327), .B2(n_0_162), 
      .ZN(n_0_161));
   INV_X1 i_0_191 (.A(n_0_163), .ZN(n_0_162));
   AOI22_X1 i_0_192 (.A1(n_0_334), .A2(n_0_164), .B1(n_0_335), .B2(n_0_212), 
      .ZN(n_0_163));
   AOI22_X1 i_0_193 (.A1(b[10]), .A2(n_0_330), .B1(b[18]), .B2(n_0_226), 
      .ZN(n_0_164));
   OAI21_X1 i_0_194 (.A(n_0_165), .B1(b[11]), .B2(n_0_356), .ZN(n_35));
   AOI21_X1 i_0_195 (.A(n_0_166), .B1(b[11]), .B2(n_0_350), .ZN(n_0_165));
   OAI221_X1 i_0_196 (.A(n_0_167), .B1(n_0_306), .B2(n_0_174), .C1(n_0_301), 
      .C2(n_0_168), .ZN(n_0_166));
   AOI22_X1 i_0_197 (.A1(n_0_352), .A2(n_0_168), .B1(n_0_353), .B2(n_0_174), 
      .ZN(n_0_167));
   AOI22_X1 i_0_198 (.A1(n_0_280), .A2(n_0_169), .B1(n_0_261), .B2(n_0_189), 
      .ZN(n_0_168));
   OAI21_X1 i_0_199 (.A(n_0_170), .B1(n_0_326), .B2(n_0_171), .ZN(n_0_169));
   NAND2_X1 i_0_200 (.A1(n_0_326), .A2(n_0_203), .ZN(n_0_170));
   INV_X1 i_0_201 (.A(n_0_172), .ZN(n_0_171));
   AOI22_X1 i_0_202 (.A1(n_0_334), .A2(n_0_173), .B1(n_0_335), .B2(n_0_225), 
      .ZN(n_0_172));
   AOI22_X1 i_0_203 (.A1(b[11]), .A2(n_0_330), .B1(b[19]), .B2(n_0_226), 
      .ZN(n_0_173));
   AOI22_X1 i_0_204 (.A1(n_0_271), .A2(n_0_175), .B1(n_0_254), .B2(n_0_183), 
      .ZN(n_0_174));
   AOI22_X1 i_0_205 (.A1(n_0_310), .A2(n_0_176), .B1(n_0_309), .B2(n_0_198), 
      .ZN(n_0_175));
   OAI21_X1 i_0_206 (.A(n_0_177), .B1(n_0_322), .B2(n_0_231), .ZN(n_0_176));
   NAND2_X1 i_0_207 (.A1(n_0_322), .A2(n_0_178), .ZN(n_0_177));
   AOI22_X1 i_0_208 (.A1(a[11]), .A2(n_0_317), .B1(a[19]), .B2(n_0_232), 
      .ZN(n_0_178));
   OAI21_X1 i_0_209 (.A(n_0_179), .B1(b[12]), .B2(n_0_356), .ZN(n_36));
   AOI21_X1 i_0_210 (.A(n_0_180), .B1(b[12]), .B2(n_0_350), .ZN(n_0_179));
   OAI221_X1 i_0_211 (.A(n_0_181), .B1(n_0_306), .B2(n_0_182), .C1(n_0_301), 
      .C2(n_0_188), .ZN(n_0_180));
   AOI22_X1 i_0_212 (.A1(n_0_352), .A2(n_0_188), .B1(n_0_353), .B2(n_0_182), 
      .ZN(n_0_181));
   AOI22_X1 i_0_213 (.A1(n_0_254), .A2(n_0_197), .B1(n_0_271), .B2(n_0_183), 
      .ZN(n_0_182));
   AOI21_X1 i_0_214 (.A(n_0_184), .B1(n_0_309), .B2(n_0_216), .ZN(n_0_183));
   NOR2_X1 i_0_215 (.A1(n_0_309), .A2(n_0_185), .ZN(n_0_184));
   OAI21_X1 i_0_216 (.A(n_0_187), .B1(n_0_323), .B2(n_0_186), .ZN(n_0_185));
   AOI22_X1 i_0_217 (.A1(a[12]), .A2(n_0_317), .B1(a[20]), .B2(n_0_232), 
      .ZN(n_0_186));
   NAND2_X1 i_0_218 (.A1(a[16]), .A2(n_0_268), .ZN(n_0_187));
   AOI22_X1 i_0_219 (.A1(n_0_261), .A2(n_0_201), .B1(n_0_280), .B2(n_0_189), 
      .ZN(n_0_188));
   AOI22_X1 i_0_220 (.A1(n_0_327), .A2(n_0_190), .B1(n_0_326), .B2(n_0_210), 
      .ZN(n_0_189));
   AOI22_X1 i_0_221 (.A1(n_0_334), .A2(n_0_191), .B1(b[16]), .B2(n_0_278), 
      .ZN(n_0_190));
   INV_X1 i_0_222 (.A(n_0_192), .ZN(n_0_191));
   AOI22_X1 i_0_223 (.A1(b[12]), .A2(n_0_330), .B1(b[20]), .B2(n_0_226), 
      .ZN(n_0_192));
   OAI21_X1 i_0_224 (.A(n_0_193), .B1(b[13]), .B2(n_0_356), .ZN(n_37));
   AOI21_X1 i_0_225 (.A(n_0_194), .B1(b[13]), .B2(n_0_350), .ZN(n_0_193));
   OAI221_X1 i_0_226 (.A(n_0_195), .B1(n_0_301), .B2(n_0_200), .C1(n_0_306), 
      .C2(n_0_196), .ZN(n_0_194));
   AOI22_X1 i_0_227 (.A1(n_0_353), .A2(n_0_196), .B1(n_0_352), .B2(n_0_200), 
      .ZN(n_0_195));
   AOI22_X1 i_0_228 (.A1(n_0_271), .A2(n_0_197), .B1(n_0_254), .B2(n_0_215), 
      .ZN(n_0_196));
   AOI22_X1 i_0_229 (.A1(n_0_310), .A2(n_0_198), .B1(n_0_309), .B2(n_0_230), 
      .ZN(n_0_197));
   AOI22_X1 i_0_230 (.A1(n_0_322), .A2(n_0_199), .B1(a[17]), .B2(n_0_268), 
      .ZN(n_0_198));
   OAI33_X1 i_0_231 (.A1(n_0_321), .A2(n_0_318), .A3(n_0_489), .B1(n_0_320), 
      .B2(n_0_318), .B3(n_0_497), .ZN(n_0_199));
   AOI22_X1 i_0_232 (.A1(n_0_261), .A2(n_0_209), .B1(n_0_280), .B2(n_0_201), 
      .ZN(n_0_200));
   INV_X1 i_0_233 (.A(n_0_202), .ZN(n_0_201));
   AOI22_X1 i_0_234 (.A1(n_0_327), .A2(n_0_203), .B1(n_0_326), .B2(n_0_224), 
      .ZN(n_0_202));
   OAI21_X1 i_0_235 (.A(n_0_205), .B1(n_0_335), .B2(n_0_204), .ZN(n_0_203));
   AOI22_X1 i_0_236 (.A1(b[13]), .A2(n_0_330), .B1(b[21]), .B2(n_0_226), 
      .ZN(n_0_204));
   NAND2_X1 i_0_237 (.A1(b[17]), .A2(n_0_278), .ZN(n_0_205));
   OAI21_X1 i_0_238 (.A(n_0_206), .B1(b[14]), .B2(n_0_356), .ZN(n_38));
   AOI221_X1 i_0_239 (.A(n_0_207), .B1(n_0_352), .B2(n_0_208), .C1(b[14]), 
      .C2(n_0_350), .ZN(n_0_206));
   OAI221_X1 i_0_240 (.A(n_0_213), .B1(n_0_306), .B2(n_0_214), .C1(n_0_301), 
      .C2(n_0_208), .ZN(n_0_207));
   AOI22_X1 i_0_241 (.A1(n_0_280), .A2(n_0_209), .B1(n_0_261), .B2(n_0_222), 
      .ZN(n_0_208));
   OAI22_X1 i_0_242 (.A1(n_0_326), .A2(n_0_210), .B1(n_0_327), .B2(n_0_241), 
      .ZN(n_0_209));
   AOI21_X1 i_0_243 (.A(n_0_211), .B1(b[18]), .B2(n_0_278), .ZN(n_0_210));
   NOR2_X1 i_0_244 (.A1(n_0_335), .A2(n_0_212), .ZN(n_0_211));
   AOI22_X1 i_0_245 (.A1(b[14]), .A2(n_0_330), .B1(b[22]), .B2(n_0_226), 
      .ZN(n_0_212));
   NAND2_X1 i_0_246 (.A1(n_0_353), .A2(n_0_214), .ZN(n_0_213));
   AOI22_X1 i_0_247 (.A1(n_0_254), .A2(n_0_229), .B1(n_0_271), .B2(n_0_215), 
      .ZN(n_0_214));
   AOI22_X1 i_0_248 (.A1(n_0_310), .A2(n_0_216), .B1(n_0_309), .B2(n_0_238), 
      .ZN(n_0_215));
   AOI22_X1 i_0_249 (.A1(n_0_322), .A2(n_0_217), .B1(a[18]), .B2(n_0_268), 
      .ZN(n_0_216));
   OAI33_X1 i_0_250 (.A1(n_0_321), .A2(n_0_318), .A3(n_0_490), .B1(n_0_320), 
      .B2(n_0_318), .B3(n_0_498), .ZN(n_0_217));
   OAI21_X1 i_0_251 (.A(n_0_218), .B1(b[15]), .B2(n_0_356), .ZN(n_39));
   AOI21_X1 i_0_252 (.A(n_0_219), .B1(b[15]), .B2(n_0_350), .ZN(n_0_218));
   OAI221_X1 i_0_253 (.A(n_0_220), .B1(n_0_306), .B2(n_0_228), .C1(n_0_301), 
      .C2(n_0_221), .ZN(n_0_219));
   AOI22_X1 i_0_254 (.A1(n_0_353), .A2(n_0_228), .B1(n_0_352), .B2(n_0_221), 
      .ZN(n_0_220));
   AOI22_X1 i_0_255 (.A1(n_0_261), .A2(n_0_240), .B1(n_0_280), .B2(n_0_222), 
      .ZN(n_0_221));
   AOI21_X1 i_0_256 (.A(n_0_223), .B1(n_0_326), .B2(n_0_250), .ZN(n_0_222));
   NOR2_X1 i_0_257 (.A1(n_0_326), .A2(n_0_224), .ZN(n_0_223));
   OAI21_X1 i_0_258 (.A(n_0_227), .B1(n_0_335), .B2(n_0_225), .ZN(n_0_224));
   AOI22_X1 i_0_259 (.A1(b[15]), .A2(n_0_330), .B1(n_0_402), .B2(n_0_226), 
      .ZN(n_0_225));
   AND2_X1 i_0_260 (.A1(n_0_333), .A2(n_0_332), .ZN(n_0_226));
   NAND2_X1 i_0_261 (.A1(b[19]), .A2(n_0_278), .ZN(n_0_227));
   AOI22_X1 i_0_262 (.A1(n_0_254), .A2(n_0_237), .B1(n_0_271), .B2(n_0_229), 
      .ZN(n_0_228));
   AOI22_X1 i_0_263 (.A1(n_0_310), .A2(n_0_230), .B1(n_0_309), .B2(n_0_246), 
      .ZN(n_0_229));
   AOI22_X1 i_0_264 (.A1(n_0_322), .A2(n_0_231), .B1(a[19]), .B2(n_0_268), 
      .ZN(n_0_230));
   OAI33_X1 i_0_265 (.A1(n_0_321), .A2(n_0_318), .A3(n_0_491), .B1(n_0_320), 
      .B2(n_0_318), .B3(n_0_405), .ZN(n_0_231));
   NOR2_X1 i_0_266 (.A1(n_0_320), .A2(n_0_318), .ZN(n_0_232));
   OAI211_X1 i_0_267 (.A(n_0_233), .B(n_0_235), .C1(b[16]), .C2(n_0_356), 
      .ZN(n_40));
   AOI21_X1 i_0_268 (.A(n_0_234), .B1(n_0_353), .B2(n_0_236), .ZN(n_0_233));
   OAI22_X1 i_0_269 (.A1(n_0_301), .A2(n_0_239), .B1(n_0_306), .B2(n_0_236), 
      .ZN(n_0_234));
   AOI22_X1 i_0_270 (.A1(b[16]), .A2(n_0_350), .B1(n_0_352), .B2(n_0_239), 
      .ZN(n_0_235));
   AOI22_X1 i_0_271 (.A1(n_0_254), .A2(n_0_245), .B1(n_0_271), .B2(n_0_237), 
      .ZN(n_0_236));
   AOI22_X1 i_0_272 (.A1(n_0_310), .A2(n_0_238), .B1(n_0_309), .B2(n_0_256), 
      .ZN(n_0_237));
   AOI22_X1 i_0_273 (.A1(a[16]), .A2(n_0_316), .B1(a[20]), .B2(n_0_268), 
      .ZN(n_0_238));
   AOI22_X1 i_0_274 (.A1(n_0_261), .A2(n_0_249), .B1(n_0_280), .B2(n_0_240), 
      .ZN(n_0_239));
   AOI22_X1 i_0_275 (.A1(n_0_327), .A2(n_0_241), .B1(n_0_326), .B2(n_0_260), 
      .ZN(n_0_240));
   AOI22_X1 i_0_276 (.A1(b[16]), .A2(n_0_329), .B1(b[20]), .B2(n_0_278), 
      .ZN(n_0_241));
   OAI211_X1 i_0_277 (.A(n_0_243), .B(n_0_242), .C1(n_0_306), .C2(n_0_244), 
      .ZN(n_41));
   AOI222_X1 i_0_278 (.A1(b[17]), .A2(n_0_350), .B1(n_0_353), .B2(n_0_244), 
      .C1(n_0_523), .C2(n_0_355), .ZN(n_0_242));
   AOI22_X1 i_0_279 (.A1(n_0_352), .A2(n_0_248), .B1(n_0_302), .B2(n_0_247), 
      .ZN(n_0_243));
   AOI22_X1 i_0_280 (.A1(n_0_271), .A2(n_0_245), .B1(n_0_255), .B2(n_0_254), 
      .ZN(n_0_244));
   AOI22_X1 i_0_281 (.A1(n_0_310), .A2(n_0_246), .B1(n_0_309), .B2(n_0_267), 
      .ZN(n_0_245));
   AOI22_X1 i_0_282 (.A1(a[17]), .A2(n_0_316), .B1(a[21]), .B2(n_0_268), 
      .ZN(n_0_246));
   INV_X1 i_0_283 (.A(n_0_248), .ZN(n_0_247));
   AOI22_X1 i_0_284 (.A1(n_0_280), .A2(n_0_249), .B1(n_0_261), .B2(n_0_259), 
      .ZN(n_0_248));
   AOI22_X1 i_0_285 (.A1(n_0_327), .A2(n_0_250), .B1(n_0_326), .B2(n_0_277), 
      .ZN(n_0_249));
   AOI22_X1 i_0_286 (.A1(b[17]), .A2(n_0_329), .B1(b[21]), .B2(n_0_278), 
      .ZN(n_0_250));
   OAI211_X1 i_0_287 (.A(n_0_252), .B(n_0_251), .C1(n_0_306), .C2(n_0_253), 
      .ZN(n_42));
   AOI222_X1 i_0_288 (.A1(b[18]), .A2(n_0_350), .B1(n_0_353), .B2(n_0_253), 
      .C1(n_0_524), .C2(n_0_355), .ZN(n_0_251));
   AOI22_X1 i_0_289 (.A1(n_0_352), .A2(n_0_258), .B1(n_0_302), .B2(n_0_257), 
      .ZN(n_0_252));
   AOI22_X1 i_0_290 (.A1(n_0_271), .A2(n_0_255), .B1(n_0_266), .B2(n_0_254), 
      .ZN(n_0_253));
   AND2_X1 i_0_291 (.A1(n_0_448), .A2(n_0_312), .ZN(n_0_254));
   OAI22_X1 i_0_292 (.A1(n_0_309), .A2(n_0_256), .B1(n_0_496), .B2(n_0_269), 
      .ZN(n_0_255));
   AOI22_X1 i_0_293 (.A1(a[18]), .A2(n_0_316), .B1(a[22]), .B2(n_0_268), 
      .ZN(n_0_256));
   INV_X1 i_0_294 (.A(n_0_258), .ZN(n_0_257));
   AOI22_X1 i_0_295 (.A1(n_0_275), .A2(n_0_261), .B1(n_0_280), .B2(n_0_259), 
      .ZN(n_0_258));
   OAI22_X1 i_0_296 (.A1(n_0_326), .A2(n_0_260), .B1(n_0_526), .B2(n_0_276), 
      .ZN(n_0_259));
   AOI22_X1 i_0_297 (.A1(b[18]), .A2(n_0_329), .B1(b[22]), .B2(n_0_278), 
      .ZN(n_0_260));
   AND2_X1 i_0_298 (.A1(n_0_448), .A2(n_0_336), .ZN(n_0_261));
   OAI21_X1 i_0_299 (.A(n_0_262), .B1(b[19]), .B2(n_0_356), .ZN(n_43));
   AOI21_X1 i_0_300 (.A(n_0_263), .B1(b[19]), .B2(n_0_350), .ZN(n_0_262));
   OAI221_X1 i_0_301 (.A(n_0_264), .B1(n_0_351), .B2(n_0_273), .C1(n_0_306), 
      .C2(n_0_265), .ZN(n_0_263));
   AOI22_X1 i_0_302 (.A1(n_0_302), .A2(n_0_273), .B1(n_0_353), .B2(n_0_265), 
      .ZN(n_0_264));
   OAI21_X1 i_0_303 (.A(n_0_270), .B1(n_0_448), .B2(n_0_266), .ZN(n_0_265));
   OAI22_X1 i_0_304 (.A1(n_0_497), .A2(n_0_269), .B1(n_0_309), .B2(n_0_267), 
      .ZN(n_0_266));
   AOI22_X1 i_0_305 (.A1(a[19]), .A2(n_0_316), .B1(n_0_404), .B2(n_0_268), 
      .ZN(n_0_267));
   NOR3_X1 i_0_306 (.A1(n_0_321), .A2(n_0_318), .A3(n_0_322), .ZN(n_0_268));
   NAND2_X1 i_0_307 (.A1(n_0_316), .A2(n_0_309), .ZN(n_0_269));
   OAI21_X1 i_0_308 (.A(n_0_272), .B1(n_0_311), .B2(n_0_286), .ZN(n_0_270));
   INV_X1 i_0_309 (.A(n_0_272), .ZN(n_0_271));
   NAND2_X1 i_0_310 (.A1(n_0_447), .A2(n_0_312), .ZN(n_0_272));
   INV_X1 i_0_311 (.A(n_0_274), .ZN(n_0_273));
   OAI21_X1 i_0_312 (.A(n_0_279), .B1(n_0_448), .B2(n_0_275), .ZN(n_0_274));
   OAI22_X1 i_0_313 (.A1(n_0_326), .A2(n_0_277), .B1(n_0_527), .B2(n_0_276), 
      .ZN(n_0_275));
   NAND2_X1 i_0_314 (.A1(n_0_329), .A2(n_0_326), .ZN(n_0_276));
   AOI22_X1 i_0_315 (.A1(n_0_402), .A2(n_0_278), .B1(b[19]), .B2(n_0_329), 
      .ZN(n_0_277));
   NOR3_X1 i_0_316 (.A1(n_0_333), .A2(n_0_331), .A3(n_0_334), .ZN(n_0_278));
   OAI21_X1 i_0_317 (.A(n_0_281), .B1(n_0_328), .B2(n_0_288), .ZN(n_0_279));
   INV_X1 i_0_318 (.A(n_0_281), .ZN(n_0_280));
   NAND2_X1 i_0_319 (.A1(n_0_447), .A2(n_0_336), .ZN(n_0_281));
   OAI211_X1 i_0_320 (.A(n_0_283), .B(n_0_282), .C1(b[20]), .C2(n_0_356), 
      .ZN(n_44));
   AOI22_X1 i_0_321 (.A1(b[20]), .A2(n_0_350), .B1(n_0_305), .B2(n_0_285), 
      .ZN(n_0_282));
   AOI21_X1 i_0_322 (.A(n_0_284), .B1(n_0_302), .B2(n_0_287), .ZN(n_0_283));
   OAI22_X1 i_0_323 (.A1(n_0_351), .A2(n_0_287), .B1(n_0_354), .B2(n_0_285), 
      .ZN(n_0_284));
   AOI221_X1 i_0_324 (.A(n_0_311), .B1(n_0_448), .B2(n_0_296), .C1(n_0_447), 
      .C2(n_0_286), .ZN(n_0_285));
   AOI22_X1 i_0_325 (.A1(a[20]), .A2(n_0_310), .B1(a[22]), .B2(n_0_309), 
      .ZN(n_0_286));
   AOI221_X1 i_0_326 (.A(n_0_328), .B1(n_0_447), .B2(n_0_288), .C1(n_0_448), 
      .C2(n_0_299), .ZN(n_0_287));
   AOI22_X1 i_0_327 (.A1(b[22]), .A2(n_0_326), .B1(b[20]), .B2(n_0_327), 
      .ZN(n_0_288));
   OAI21_X1 i_0_328 (.A(n_0_289), .B1(b[21]), .B2(n_0_356), .ZN(n_45));
   AOI21_X1 i_0_329 (.A(n_0_290), .B1(b[21]), .B2(n_0_350), .ZN(n_0_289));
   OAI21_X1 i_0_330 (.A(n_0_291), .B1(n_0_351), .B2(n_0_297), .ZN(n_0_290));
   AOI21_X1 i_0_331 (.A(n_0_292), .B1(n_0_302), .B2(n_0_297), .ZN(n_0_291));
   AOI22_X1 i_0_332 (.A1(n_0_354), .A2(n_0_293), .B1(n_0_306), .B2(n_0_294), 
      .ZN(n_0_292));
   INV_X1 i_0_333 (.A(n_0_294), .ZN(n_0_293));
   AOI211_X1 i_0_334 (.A(n_0_295), .B(n_0_311), .C1(n_0_447), .C2(n_0_296), 
      .ZN(n_0_294));
   AOI21_X1 i_0_335 (.A(n_0_447), .B1(a[22]), .B2(n_0_310), .ZN(n_0_295));
   OAI22_X1 i_0_336 (.A1(a[21]), .A2(n_0_309), .B1(n_0_404), .B2(n_0_310), 
      .ZN(n_0_296));
   AOI211_X1 i_0_337 (.A(n_0_298), .B(n_0_328), .C1(n_0_447), .C2(n_0_299), 
      .ZN(n_0_297));
   AOI21_X1 i_0_338 (.A(n_0_447), .B1(b[22]), .B2(n_0_327), .ZN(n_0_298));
   AOI22_X1 i_0_339 (.A1(n_0_402), .A2(n_0_326), .B1(b[21]), .B2(n_0_327), 
      .ZN(n_0_299));
   OAI211_X1 i_0_340 (.A(n_0_300), .B(n_0_303), .C1(b[22]), .C2(n_0_356), 
      .ZN(n_46));
   AOI22_X1 i_0_341 (.A1(b[22]), .A2(n_0_350), .B1(n_0_324), .B2(n_0_302), 
      .ZN(n_0_300));
   INV_X1 i_0_342 (.A(n_0_302), .ZN(n_0_301));
   NOR2_X1 i_0_343 (.A1(n_0_450), .A2(n_0_398), .ZN(n_0_302));
   AOI21_X1 i_0_344 (.A(n_0_304), .B1(n_0_307), .B2(n_0_305), .ZN(n_0_303));
   OAI22_X1 i_0_345 (.A1(n_0_351), .A2(n_0_324), .B1(n_0_354), .B2(n_0_307), 
      .ZN(n_0_304));
   INV_X1 i_0_346 (.A(n_0_306), .ZN(n_0_305));
   NAND2_X1 i_0_347 (.A1(n_0_437), .A2(n_0_399), .ZN(n_0_306));
   AOI211_X1 i_0_348 (.A(n_0_311), .B(n_0_308), .C1(n_0_498), .C2(n_0_447), 
      .ZN(n_0_307));
   OAI21_X1 i_0_349 (.A(n_0_310), .B1(n_0_466), .B2(n_0_404), .ZN(n_0_308));
   INV_X1 i_0_350 (.A(n_0_310), .ZN(n_0_309));
   XNOR2_X1 i_0_351 (.A(n_0_465), .B(n_0_464), .ZN(n_0_310));
   NAND2_X1 i_0_352 (.A1(n_0_316), .A2(n_0_312), .ZN(n_0_311));
   AOI221_X1 i_0_353 (.A(n_0_313), .B1(n_0_476), .B2(n_0_442), .C1(n_0_454), 
      .C2(n_0_315), .ZN(n_0_312));
   AOI22_X1 i_0_354 (.A1(n_0_456), .A2(n_0_314), .B1(n_0_474), .B2(n_0_315), 
      .ZN(n_0_313));
   OAI22_X1 i_0_355 (.A1(b[28]), .A2(n_0_504), .B1(n_0_452), .B2(n_0_442), 
      .ZN(n_0_314));
   NOR2_X1 i_0_356 (.A1(n_0_452), .A2(n_0_442), .ZN(n_0_315));
   NOR3_X1 i_0_357 (.A1(n_0_321), .A2(n_0_318), .A3(n_0_323), .ZN(n_0_316));
   NOR2_X1 i_0_358 (.A1(n_0_321), .A2(n_0_318), .ZN(n_0_317));
   INV_X1 i_0_359 (.A(n_0_319), .ZN(n_0_318));
   XNOR2_X1 i_0_360 (.A(n_0_459), .B(n_0_458), .ZN(n_0_319));
   INV_X1 i_0_361 (.A(n_0_321), .ZN(n_0_320));
   XNOR2_X1 i_0_362 (.A(n_0_473), .B(n_0_460), .ZN(n_0_321));
   INV_X1 i_0_363 (.A(n_0_323), .ZN(n_0_322));
   OAI21_X1 i_0_364 (.A(n_0_461), .B1(n_0_472), .B2(n_0_462), .ZN(n_0_323));
   AOI211_X1 i_0_365 (.A(n_0_328), .B(n_0_325), .C1(n_0_528), .C2(n_0_447), 
      .ZN(n_0_324));
   OAI21_X1 i_0_366 (.A(n_0_327), .B1(n_0_469), .B2(n_0_402), .ZN(n_0_325));
   INV_X1 i_0_367 (.A(n_0_327), .ZN(n_0_326));
   XNOR2_X1 i_0_368 (.A(n_0_464), .B(n_0_449), .ZN(n_0_327));
   NAND2_X1 i_0_369 (.A1(n_0_336), .A2(n_0_329), .ZN(n_0_328));
   NOR3_X1 i_0_370 (.A1(n_0_333), .A2(n_0_331), .A3(n_0_335), .ZN(n_0_329));
   NOR2_X1 i_0_371 (.A1(n_0_333), .A2(n_0_331), .ZN(n_0_330));
   INV_X1 i_0_372 (.A(n_0_332), .ZN(n_0_331));
   XNOR2_X1 i_0_373 (.A(n_0_457), .B(n_0_344), .ZN(n_0_332));
   OAI21_X1 i_0_374 (.A(n_0_345), .B1(n_0_473), .B2(n_0_346), .ZN(n_0_333));
   INV_X1 i_0_375 (.A(n_0_335), .ZN(n_0_334));
   OAI21_X1 i_0_376 (.A(n_0_347), .B1(n_0_472), .B2(n_0_348), .ZN(n_0_335));
   AOI21_X1 i_0_377 (.A(n_0_337), .B1(n_0_442), .B2(n_0_341), .ZN(n_0_336));
   OAI21_X1 i_0_378 (.A(n_0_338), .B1(n_0_442), .B2(n_0_341), .ZN(n_0_337));
   OAI21_X1 i_0_379 (.A(n_0_342), .B1(n_0_445), .B2(n_0_339), .ZN(n_0_338));
   INV_X1 i_0_380 (.A(n_0_340), .ZN(n_0_339));
   AOI21_X1 i_0_381 (.A(n_0_343), .B1(n_0_474), .B2(n_0_446), .ZN(n_0_340));
   AOI21_X1 i_0_382 (.A(n_0_452), .B1(n_0_475), .B2(n_0_342), .ZN(n_0_341));
   NAND2_X1 i_0_383 (.A1(n_0_444), .A2(n_0_343), .ZN(n_0_342));
   AOI22_X1 i_0_384 (.A1(b[27]), .A2(n_0_503), .B1(n_0_458), .B2(n_0_344), 
      .ZN(n_0_343));
   OAI21_X1 i_0_385 (.A(n_0_345), .B1(n_0_532), .B2(a[26]), .ZN(n_0_344));
   NAND2_X1 i_0_386 (.A1(n_0_473), .A2(n_0_346), .ZN(n_0_345));
   OAI21_X1 i_0_387 (.A(n_0_347), .B1(n_0_531), .B2(a[25]), .ZN(n_0_346));
   NAND2_X1 i_0_388 (.A1(n_0_472), .A2(n_0_348), .ZN(n_0_347));
   OAI22_X1 i_0_389 (.A1(n_0_530), .A2(a[24]), .B1(n_0_463), .B2(n_0_449), 
      .ZN(n_0_348));
   OAI21_X1 i_0_390 (.A(n_0_349), .B1(n_0_402), .B2(n_0_356), .ZN(n_47));
   AOI211_X1 i_0_391 (.A(n_0_353), .B(n_0_352), .C1(n_0_402), .C2(n_0_350), 
      .ZN(n_0_349));
   NOR2_X1 i_0_392 (.A1(n_0_440), .A2(n_0_357), .ZN(n_0_350));
   INV_X1 i_0_393 (.A(n_0_352), .ZN(n_0_351));
   NOR2_X1 i_0_394 (.A1(n_0_450), .A2(n_0_399), .ZN(n_0_352));
   INV_X1 i_0_395 (.A(n_0_354), .ZN(n_0_353));
   NAND2_X1 i_0_396 (.A1(n_0_437), .A2(n_0_398), .ZN(n_0_354));
   INV_X1 i_0_397 (.A(n_0_356), .ZN(n_0_355));
   NAND2_X1 i_0_398 (.A1(n_0_439), .A2(n_0_357), .ZN(n_0_356));
   NOR2_X1 i_0_399 (.A1(n_0_400), .A2(n_0_399), .ZN(n_0_357));
   INV_X1 i_0_400 (.A(n_0_358), .ZN(out[0]));
   AOI22_X1 i_0_401 (.A1(CLA_SUM[0]), .A2(n_0_389), .B1(CLA_SUM[1]), .B2(n_0_391), 
      .ZN(n_0_358));
   INV_X1 i_0_402 (.A(n_0_359), .ZN(out[1]));
   AOI222_X1 i_0_403 (.A1(o_m[1]), .A2(n_48), .B1(CLA_SUM[2]), .B2(n_0_391), 
      .C1(CLA_SUM[1]), .C2(n_0_389), .ZN(n_0_359));
   INV_X1 i_0_404 (.A(n_0_360), .ZN(out[2]));
   AOI222_X1 i_0_405 (.A1(o_m[2]), .A2(n_48), .B1(CLA_SUM[3]), .B2(n_0_391), 
      .C1(CLA_SUM[2]), .C2(n_0_389), .ZN(n_0_360));
   INV_X1 i_0_406 (.A(n_0_361), .ZN(out[3]));
   AOI222_X1 i_0_407 (.A1(o_m[3]), .A2(n_48), .B1(CLA_SUM[4]), .B2(n_0_391), 
      .C1(CLA_SUM[3]), .C2(n_0_389), .ZN(n_0_361));
   INV_X1 i_0_408 (.A(n_0_362), .ZN(out[4]));
   AOI222_X1 i_0_409 (.A1(o_m[4]), .A2(n_48), .B1(CLA_SUM[5]), .B2(n_0_391), 
      .C1(CLA_SUM[4]), .C2(n_0_389), .ZN(n_0_362));
   INV_X1 i_0_410 (.A(n_0_363), .ZN(out[5]));
   AOI222_X1 i_0_411 (.A1(o_m[5]), .A2(n_48), .B1(CLA_SUM[6]), .B2(n_0_391), 
      .C1(CLA_SUM[5]), .C2(n_0_389), .ZN(n_0_363));
   INV_X1 i_0_412 (.A(n_0_364), .ZN(out[6]));
   AOI222_X1 i_0_413 (.A1(o_m[6]), .A2(n_48), .B1(CLA_SUM[7]), .B2(n_0_391), 
      .C1(CLA_SUM[6]), .C2(n_0_389), .ZN(n_0_364));
   INV_X1 i_0_414 (.A(n_0_365), .ZN(out[7]));
   AOI222_X1 i_0_415 (.A1(o_m[7]), .A2(n_48), .B1(CLA_SUM[8]), .B2(n_0_391), 
      .C1(CLA_SUM[7]), .C2(n_0_389), .ZN(n_0_365));
   INV_X1 i_0_416 (.A(n_0_366), .ZN(out[8]));
   AOI222_X1 i_0_417 (.A1(o_m[8]), .A2(n_48), .B1(CLA_SUM[9]), .B2(n_0_391), 
      .C1(CLA_SUM[8]), .C2(n_0_389), .ZN(n_0_366));
   INV_X1 i_0_418 (.A(n_0_367), .ZN(out[9]));
   AOI222_X1 i_0_419 (.A1(o_m[9]), .A2(n_48), .B1(CLA_SUM[10]), .B2(n_0_391), 
      .C1(CLA_SUM[9]), .C2(n_0_389), .ZN(n_0_367));
   INV_X1 i_0_420 (.A(n_0_368), .ZN(out[10]));
   AOI222_X1 i_0_421 (.A1(o_m[10]), .A2(n_48), .B1(CLA_SUM[11]), .B2(n_0_391), 
      .C1(CLA_SUM[10]), .C2(n_0_389), .ZN(n_0_368));
   INV_X1 i_0_422 (.A(n_0_369), .ZN(out[11]));
   AOI222_X1 i_0_423 (.A1(o_m[11]), .A2(n_48), .B1(CLA_SUM[12]), .B2(n_0_391), 
      .C1(CLA_SUM[11]), .C2(n_0_389), .ZN(n_0_369));
   INV_X1 i_0_424 (.A(n_0_370), .ZN(out[12]));
   AOI222_X1 i_0_425 (.A1(o_m[12]), .A2(n_48), .B1(CLA_SUM[13]), .B2(n_0_391), 
      .C1(CLA_SUM[12]), .C2(n_0_389), .ZN(n_0_370));
   INV_X1 i_0_426 (.A(n_0_371), .ZN(out[13]));
   AOI222_X1 i_0_427 (.A1(o_m[13]), .A2(n_48), .B1(CLA_SUM[14]), .B2(n_0_391), 
      .C1(CLA_SUM[13]), .C2(n_0_389), .ZN(n_0_371));
   INV_X1 i_0_428 (.A(n_0_372), .ZN(out[14]));
   AOI222_X1 i_0_429 (.A1(o_m[14]), .A2(n_48), .B1(CLA_SUM[15]), .B2(n_0_391), 
      .C1(CLA_SUM[14]), .C2(n_0_389), .ZN(n_0_372));
   INV_X1 i_0_430 (.A(n_0_373), .ZN(out[15]));
   AOI222_X1 i_0_431 (.A1(o_m[15]), .A2(n_48), .B1(CLA_SUM[16]), .B2(n_0_391), 
      .C1(CLA_SUM[15]), .C2(n_0_389), .ZN(n_0_373));
   INV_X1 i_0_432 (.A(n_0_374), .ZN(out[16]));
   AOI222_X1 i_0_433 (.A1(o_m[16]), .A2(n_48), .B1(CLA_SUM[17]), .B2(n_0_391), 
      .C1(CLA_SUM[16]), .C2(n_0_389), .ZN(n_0_374));
   INV_X1 i_0_434 (.A(n_0_375), .ZN(out[17]));
   AOI222_X1 i_0_435 (.A1(o_m[17]), .A2(n_48), .B1(CLA_SUM[18]), .B2(n_0_391), 
      .C1(CLA_SUM[17]), .C2(n_0_389), .ZN(n_0_375));
   INV_X1 i_0_436 (.A(n_0_376), .ZN(out[18]));
   AOI222_X1 i_0_437 (.A1(o_m[18]), .A2(n_48), .B1(CLA_SUM[19]), .B2(n_0_391), 
      .C1(CLA_SUM[18]), .C2(n_0_389), .ZN(n_0_376));
   INV_X1 i_0_438 (.A(n_0_377), .ZN(out[19]));
   AOI222_X1 i_0_439 (.A1(o_m[19]), .A2(n_48), .B1(CLA_SUM[20]), .B2(n_0_391), 
      .C1(CLA_SUM[19]), .C2(n_0_389), .ZN(n_0_377));
   INV_X1 i_0_440 (.A(n_0_378), .ZN(out[20]));
   AOI222_X1 i_0_441 (.A1(o_m[20]), .A2(n_48), .B1(CLA_SUM[21]), .B2(n_0_391), 
      .C1(CLA_SUM[20]), .C2(n_0_389), .ZN(n_0_378));
   INV_X1 i_0_442 (.A(n_0_379), .ZN(out[21]));
   AOI222_X1 i_0_443 (.A1(o_m[21]), .A2(n_48), .B1(CLA_SUM[22]), .B2(n_0_391), 
      .C1(CLA_SUM[21]), .C2(n_0_389), .ZN(n_0_379));
   AOI21_X1 i_0_444 (.A(n_0_380), .B1(n_0_479), .B2(n_0_389), .ZN(out[22]));
   AOI21_X1 i_0_445 (.A(CLA_SUM[23]), .B1(o_m[22]), .B2(n_0_392), .ZN(n_0_380));
   OAI21_X1 i_0_446 (.A(n_0_381), .B1(n_49), .B2(n_0_392), .ZN(out[23]));
   AOI22_X1 i_0_447 (.A1(o_e[0]), .A2(n_48), .B1(n_49), .B2(n_0_389), .ZN(
      n_0_381));
   INV_X1 i_0_448 (.A(n_0_382), .ZN(out[24]));
   AOI222_X1 i_0_449 (.A1(o_e[1]), .A2(n_48), .B1(n_0_6), .B2(n_0_391), .C1(n_50), 
      .C2(n_0_389), .ZN(n_0_382));
   INV_X1 i_0_450 (.A(n_0_383), .ZN(out[25]));
   AOI222_X1 i_0_451 (.A1(o_e[2]), .A2(n_48), .B1(n_0_7), .B2(n_0_391), .C1(n_51), 
      .C2(n_0_389), .ZN(n_0_383));
   INV_X1 i_0_452 (.A(n_0_384), .ZN(out[26]));
   AOI222_X1 i_0_453 (.A1(o_e[3]), .A2(n_48), .B1(n_0_8), .B2(n_0_391), .C1(n_52), 
      .C2(n_0_389), .ZN(n_0_384));
   INV_X1 i_0_454 (.A(n_0_385), .ZN(out[27]));
   AOI222_X1 i_0_455 (.A1(n_0_9), .A2(n_0_391), .B1(o_e[4]), .B2(n_48), .C1(n_53), 
      .C2(n_0_389), .ZN(n_0_385));
   INV_X1 i_0_456 (.A(n_0_386), .ZN(out[28]));
   AOI222_X1 i_0_457 (.A1(o_e[5]), .A2(n_48), .B1(n_0_10), .B2(n_0_391), 
      .C1(n_54), .C2(n_0_389), .ZN(n_0_386));
   INV_X1 i_0_458 (.A(n_0_387), .ZN(out[29]));
   AOI222_X1 i_0_459 (.A1(o_e[6]), .A2(n_48), .B1(n_0_11), .B2(n_0_391), 
      .C1(n_55), .C2(n_0_389), .ZN(n_0_387));
   INV_X1 i_0_460 (.A(n_0_388), .ZN(out[30]));
   AOI221_X1 i_0_461 (.A(n_0_390), .B1(o_e[7]), .B2(n_48), .C1(n_56), .C2(
      n_0_389), .ZN(n_0_388));
   AND2_X1 i_0_462 (.A1(CLA_SUM[23]), .A2(n_0_392), .ZN(n_0_389));
   AOI221_X1 i_0_463 (.A(n_0_392), .B1(n_0_478), .B2(n_0_477), .C1(n_0_5), 
      .C2(n_56), .ZN(n_0_390));
   NOR2_X1 i_0_464 (.A1(CLA_SUM[23]), .A2(n_0_391), .ZN(n_48));
   INV_X1 i_0_465 (.A(n_0_392), .ZN(n_0_391));
   OAI21_X1 i_0_466 (.A(n_0_399), .B1(CLA_COUT), .B2(n_0_439), .ZN(n_0_392));
   INV_X1 i_0_467 (.A(n_0_393), .ZN(out[31]));
   AOI22_X1 i_0_468 (.A1(a[31]), .A2(n_0_394), .B1(b[31]), .B2(n_0_395), 
      .ZN(n_0_393));
   INV_X1 i_0_469 (.A(n_0_395), .ZN(n_0_394));
   NAND2_X1 i_0_470 (.A1(n_0_438), .A2(n_0_397), .ZN(n_0_395));
   INV_X1 i_0_471 (.A(n_0_397), .ZN(n_0_396));
   NAND3_X1 i_0_472 (.A1(n_0_439), .A2(n_0_398), .A3(n_0_400), .ZN(n_0_397));
   INV_X1 i_0_473 (.A(n_0_399), .ZN(n_0_398));
   XNOR2_X1 i_0_474 (.A(b[31]), .B(a[31]), .ZN(n_0_399));
   AOI22_X1 i_0_475 (.A1(n_0_406), .A2(n_0_401), .B1(n_0_404), .B2(n_0_403), 
      .ZN(n_0_400));
   AOI22_X1 i_0_476 (.A1(n_0_405), .A2(n_0_402), .B1(b[22]), .B2(n_0_498), 
      .ZN(n_0_401));
   INV_X1 i_0_477 (.A(n_0_403), .ZN(n_0_402));
   NOR2_X1 i_0_478 (.A1(b[23]), .A2(n_0_467), .ZN(n_0_403));
   INV_X1 i_0_479 (.A(n_0_405), .ZN(n_0_404));
   NOR2_X1 i_0_480 (.A1(a[23]), .A2(n_0_470), .ZN(n_0_405));
   INV_X1 i_0_481 (.A(n_0_407), .ZN(n_0_406));
   AOI221_X1 i_0_482 (.A(n_0_408), .B1(n_0_527), .B2(a[21]), .C1(n_0_528), 
      .C2(a[22]), .ZN(n_0_407));
   AOI221_X1 i_0_483 (.A(n_0_409), .B1(b[20]), .B2(n_0_496), .C1(b[21]), 
      .C2(n_0_497), .ZN(n_0_408));
   AOI222_X1 i_0_484 (.A1(n_0_526), .A2(a[20]), .B1(n_0_525), .B2(a[19]), 
      .C1(n_0_412), .C2(n_0_410), .ZN(n_0_409));
   AOI221_X1 i_0_485 (.A(n_0_411), .B1(b[19]), .B2(n_0_495), .C1(b[18]), 
      .C2(n_0_494), .ZN(n_0_410));
   AOI211_X1 i_0_486 (.A(n_0_523), .B(a[17]), .C1(n_0_524), .C2(a[18]), .ZN(
      n_0_411));
   OAI221_X1 i_0_487 (.A(n_0_413), .B1(b[16]), .B2(n_0_492), .C1(b[17]), 
      .C2(n_0_493), .ZN(n_0_412));
   AOI21_X1 i_0_488 (.A(n_0_414), .B1(n_0_524), .B2(a[18]), .ZN(n_0_413));
   AOI21_X1 i_0_489 (.A(n_0_415), .B1(b[16]), .B2(n_0_492), .ZN(n_0_414));
   AOI22_X1 i_0_490 (.A1(n_0_522), .A2(a[15]), .B1(n_0_418), .B2(n_0_416), 
      .ZN(n_0_415));
   AOI221_X1 i_0_491 (.A(n_0_417), .B1(b[15]), .B2(n_0_491), .C1(b[14]), 
      .C2(n_0_490), .ZN(n_0_416));
   AOI211_X1 i_0_492 (.A(n_0_520), .B(a[13]), .C1(n_0_521), .C2(a[14]), .ZN(
      n_0_417));
   OAI221_X1 i_0_493 (.A(n_0_419), .B1(b[13]), .B2(n_0_489), .C1(b[14]), 
      .C2(n_0_490), .ZN(n_0_418));
   AOI21_X1 i_0_494 (.A(n_0_420), .B1(n_0_519), .B2(a[12]), .ZN(n_0_419));
   AOI21_X1 i_0_495 (.A(n_0_421), .B1(b[12]), .B2(n_0_488), .ZN(n_0_420));
   AOI22_X1 i_0_496 (.A1(n_0_423), .A2(n_0_422), .B1(n_0_518), .B2(a[11]), 
      .ZN(n_0_421));
   AOI22_X1 i_0_497 (.A1(b[11]), .A2(n_0_487), .B1(b[10]), .B2(n_0_486), 
      .ZN(n_0_422));
   INV_X1 i_0_498 (.A(n_0_424), .ZN(n_0_423));
   AOI221_X1 i_0_499 (.A(n_0_425), .B1(n_0_516), .B2(a[9]), .C1(n_0_517), 
      .C2(a[10]), .ZN(n_0_424));
   AOI221_X1 i_0_500 (.A(n_0_426), .B1(b[9]), .B2(n_0_485), .C1(b[8]), .C2(
      n_0_484), .ZN(n_0_425));
   AOI222_X1 i_0_501 (.A1(n_0_514), .A2(a[7]), .B1(n_0_515), .B2(a[8]), .C1(
      n_0_429), .C2(n_0_427), .ZN(n_0_426));
   AOI221_X1 i_0_502 (.A(n_0_428), .B1(b[7]), .B2(n_0_483), .C1(b[6]), .C2(
      n_0_482), .ZN(n_0_427));
   AOI211_X1 i_0_503 (.A(n_0_512), .B(a[5]), .C1(n_0_513), .C2(a[6]), .ZN(
      n_0_428));
   OAI221_X1 i_0_504 (.A(n_0_430), .B1(n_0_432), .B2(n_0_431), .C1(b[4]), 
      .C2(n_0_481), .ZN(n_0_429));
   AOI22_X1 i_0_505 (.A1(n_0_512), .A2(a[5]), .B1(n_0_513), .B2(a[6]), .ZN(
      n_0_430));
   OAI22_X1 i_0_506 (.A1(n_0_510), .A2(a[3]), .B1(n_0_511), .B2(a[4]), .ZN(
      n_0_431));
   AOI21_X1 i_0_507 (.A(n_0_433), .B1(n_0_510), .B2(a[3]), .ZN(n_0_432));
   AOI22_X1 i_0_508 (.A1(b[2]), .A2(n_0_480), .B1(n_0_435), .B2(n_0_434), 
      .ZN(n_0_433));
   AOI22_X1 i_0_509 (.A1(n_0_509), .A2(a[2]), .B1(n_0_508), .B2(a[1]), .ZN(
      n_0_434));
   OAI211_X1 i_0_510 (.A(n_0_507), .B(a[0]), .C1(n_0_508), .C2(a[1]), .ZN(
      n_0_435));
   INV_X1 i_0_511 (.A(n_0_436), .ZN(n_49));
   AOI22_X1 i_0_512 (.A1(n_0_466), .A2(n_0_437), .B1(n_0_469), .B2(n_0_438), 
      .ZN(n_0_436));
   AOI22_X1 i_0_513 (.A1(n_0_530), .A2(n_0_437), .B1(n_0_500), .B2(n_0_438), 
      .ZN(n_50));
   OAI22_X1 i_0_514 (.A1(n_0_531), .A2(n_0_438), .B1(n_0_501), .B2(n_0_437), 
      .ZN(n_51));
   OAI22_X1 i_0_515 (.A1(n_0_532), .A2(n_0_438), .B1(n_0_502), .B2(n_0_437), 
      .ZN(n_52));
   AOI22_X1 i_0_516 (.A1(n_0_503), .A2(n_0_438), .B1(n_0_533), .B2(n_0_437), 
      .ZN(n_53));
   AOI22_X1 i_0_517 (.A1(n_0_534), .A2(n_0_437), .B1(n_0_504), .B2(n_0_438), 
      .ZN(n_54));
   OAI22_X1 i_0_518 (.A1(n_0_535), .A2(n_0_438), .B1(n_0_505), .B2(n_0_437), 
      .ZN(n_55));
   INV_X1 i_0_519 (.A(n_0_438), .ZN(n_0_437));
   NAND2_X1 i_0_520 (.A1(n_0_450), .A2(n_0_440), .ZN(n_0_438));
   INV_X1 i_0_521 (.A(n_0_440), .ZN(n_0_439));
   NAND4_X1 i_0_522 (.A1(n_0_447), .A2(n_0_441), .A3(n_0_444), .A4(n_0_443), 
      .ZN(n_0_440));
   AND4_X1 i_0_523 (.A1(n_0_473), .A2(n_0_472), .A3(n_0_458), .A4(n_0_464), 
      .ZN(n_0_441));
   INV_X1 i_0_524 (.A(n_0_443), .ZN(n_0_442));
   AOI22_X1 i_0_525 (.A1(n_0_536), .A2(a[30]), .B1(b[30]), .B2(n_0_506), 
      .ZN(n_0_443));
   AND2_X1 i_0_526 (.A1(n_0_474), .A2(n_0_445), .ZN(n_0_444));
   AND2_X1 i_0_527 (.A1(n_0_475), .A2(n_0_453), .ZN(n_0_445));
   NAND2_X1 i_0_528 (.A1(n_0_476), .A2(n_0_453), .ZN(n_0_446));
   INV_X1 i_0_529 (.A(n_0_448), .ZN(n_0_447));
   NAND2_X1 i_0_530 (.A1(n_0_465), .A2(n_0_449), .ZN(n_0_448));
   NAND3_X1 i_0_531 (.A1(n_0_499), .A2(n_0_470), .A3(n_0_466), .ZN(n_0_449));
   AOI22_X1 i_0_532 (.A1(n_0_536), .A2(a[30]), .B1(n_0_454), .B2(n_0_451), 
      .ZN(n_0_450));
   AOI21_X1 i_0_533 (.A(n_0_452), .B1(b[30]), .B2(n_0_506), .ZN(n_0_451));
   INV_X1 i_0_534 (.A(n_0_453), .ZN(n_0_452));
   NAND2_X1 i_0_535 (.A1(b[29]), .A2(n_0_505), .ZN(n_0_453));
   NAND2_X1 i_0_536 (.A1(n_0_475), .A2(n_0_455), .ZN(n_0_454));
   NAND2_X1 i_0_537 (.A1(n_0_474), .A2(n_0_456), .ZN(n_0_455));
   OAI22_X1 i_0_538 (.A1(b[27]), .A2(n_0_503), .B1(n_0_459), .B2(n_0_457), 
      .ZN(n_0_456));
   INV_X1 i_0_539 (.A(n_0_458), .ZN(n_0_457));
   AOI22_X1 i_0_540 (.A1(n_0_533), .A2(a[27]), .B1(b[27]), .B2(n_0_503), 
      .ZN(n_0_458));
   AOI22_X1 i_0_541 (.A1(n_0_532), .A2(a[26]), .B1(n_0_473), .B2(n_0_460), 
      .ZN(n_0_459));
   OAI21_X1 i_0_542 (.A(n_0_461), .B1(b[25]), .B2(n_0_501), .ZN(n_0_460));
   NAND2_X1 i_0_543 (.A1(n_0_472), .A2(n_0_462), .ZN(n_0_461));
   OAI22_X1 i_0_544 (.A1(b[24]), .A2(n_0_500), .B1(n_0_465), .B2(n_0_463), 
      .ZN(n_0_462));
   INV_X1 i_0_545 (.A(n_0_464), .ZN(n_0_463));
   AOI22_X1 i_0_546 (.A1(n_0_530), .A2(a[24]), .B1(b[24]), .B2(n_0_500), 
      .ZN(n_0_464));
   NAND3_X1 i_0_547 (.A1(n_0_529), .A2(n_0_467), .A3(n_0_469), .ZN(n_0_465));
   NAND2_X1 i_0_548 (.A1(n_0_529), .A2(n_0_467), .ZN(n_0_466));
   NAND4_X1 i_0_549 (.A1(n_0_535), .A2(n_0_534), .A3(n_0_531), .A4(n_0_468), 
      .ZN(n_0_467));
   NOR4_X1 i_0_550 (.A1(b[30]), .A2(b[27]), .A3(b[26]), .A4(b[24]), .ZN(n_0_468));
   NAND2_X1 i_0_551 (.A1(n_0_499), .A2(n_0_470), .ZN(n_0_469));
   NAND4_X1 i_0_552 (.A1(n_0_505), .A2(n_0_504), .A3(n_0_501), .A4(n_0_471), 
      .ZN(n_0_470));
   NOR4_X1 i_0_553 (.A1(a[26]), .A2(a[24]), .A3(a[30]), .A4(a[27]), .ZN(n_0_471));
   AOI22_X1 i_0_554 (.A1(n_0_531), .A2(a[25]), .B1(b[25]), .B2(n_0_501), 
      .ZN(n_0_472));
   AOI22_X1 i_0_555 (.A1(n_0_532), .A2(a[26]), .B1(b[26]), .B2(n_0_502), 
      .ZN(n_0_473));
   NAND2_X1 i_0_556 (.A1(b[28]), .A2(n_0_504), .ZN(n_0_474));
   AOI22_X1 i_0_557 (.A1(n_0_535), .A2(a[29]), .B1(n_0_534), .B2(a[28]), 
      .ZN(n_0_475));
   NAND2_X1 i_0_558 (.A1(n_0_535), .A2(a[29]), .ZN(n_0_476));
   INV_X1 i_0_559 (.A(n_56), .ZN(n_0_477));
   NAND2_X1 i_0_560 (.A1(n_0_536), .A2(n_0_506), .ZN(n_56));
   INV_X1 i_0_561 (.A(n_0_5), .ZN(n_0_478));
   INV_X1 i_0_562 (.A(CLA_SUM[22]), .ZN(n_0_479));
   INV_X1 i_0_563 (.A(a[2]), .ZN(n_0_480));
   INV_X1 i_0_564 (.A(a[4]), .ZN(n_0_481));
   INV_X1 i_0_565 (.A(a[6]), .ZN(n_0_482));
   INV_X1 i_0_566 (.A(a[7]), .ZN(n_0_483));
   INV_X1 i_0_567 (.A(a[8]), .ZN(n_0_484));
   INV_X1 i_0_568 (.A(a[9]), .ZN(n_0_485));
   INV_X1 i_0_569 (.A(a[10]), .ZN(n_0_486));
   INV_X1 i_0_570 (.A(a[11]), .ZN(n_0_487));
   INV_X1 i_0_571 (.A(a[12]), .ZN(n_0_488));
   INV_X1 i_0_572 (.A(a[13]), .ZN(n_0_489));
   INV_X1 i_0_573 (.A(a[14]), .ZN(n_0_490));
   INV_X1 i_0_574 (.A(a[15]), .ZN(n_0_491));
   INV_X1 i_0_575 (.A(a[16]), .ZN(n_0_492));
   INV_X1 i_0_576 (.A(a[17]), .ZN(n_0_493));
   INV_X1 i_0_577 (.A(a[18]), .ZN(n_0_494));
   INV_X1 i_0_578 (.A(a[19]), .ZN(n_0_495));
   INV_X1 i_0_579 (.A(a[20]), .ZN(n_0_496));
   INV_X1 i_0_580 (.A(a[21]), .ZN(n_0_497));
   INV_X1 i_0_581 (.A(a[22]), .ZN(n_0_498));
   INV_X1 i_0_582 (.A(a[23]), .ZN(n_0_499));
   INV_X1 i_0_583 (.A(a[24]), .ZN(n_0_500));
   INV_X1 i_0_584 (.A(a[25]), .ZN(n_0_501));
   INV_X1 i_0_585 (.A(a[26]), .ZN(n_0_502));
   INV_X1 i_0_586 (.A(a[27]), .ZN(n_0_503));
   INV_X1 i_0_587 (.A(a[28]), .ZN(n_0_504));
   INV_X1 i_0_588 (.A(a[29]), .ZN(n_0_505));
   INV_X1 i_0_589 (.A(a[30]), .ZN(n_0_506));
   INV_X1 i_0_590 (.A(b[0]), .ZN(n_0_507));
   INV_X1 i_0_591 (.A(b[1]), .ZN(n_0_508));
   INV_X1 i_0_592 (.A(b[2]), .ZN(n_0_509));
   INV_X1 i_0_593 (.A(b[3]), .ZN(n_0_510));
   INV_X1 i_0_594 (.A(b[4]), .ZN(n_0_511));
   INV_X1 i_0_595 (.A(b[5]), .ZN(n_0_512));
   INV_X1 i_0_596 (.A(b[6]), .ZN(n_0_513));
   INV_X1 i_0_597 (.A(b[7]), .ZN(n_0_514));
   INV_X1 i_0_598 (.A(b[8]), .ZN(n_0_515));
   INV_X1 i_0_599 (.A(b[9]), .ZN(n_0_516));
   INV_X1 i_0_600 (.A(b[10]), .ZN(n_0_517));
   INV_X1 i_0_601 (.A(b[11]), .ZN(n_0_518));
   INV_X1 i_0_602 (.A(b[12]), .ZN(n_0_519));
   INV_X1 i_0_603 (.A(b[13]), .ZN(n_0_520));
   INV_X1 i_0_604 (.A(b[14]), .ZN(n_0_521));
   INV_X1 i_0_605 (.A(b[15]), .ZN(n_0_522));
   INV_X1 i_0_606 (.A(b[17]), .ZN(n_0_523));
   INV_X1 i_0_607 (.A(b[18]), .ZN(n_0_524));
   INV_X1 i_0_608 (.A(b[19]), .ZN(n_0_525));
   INV_X1 i_0_609 (.A(b[20]), .ZN(n_0_526));
   INV_X1 i_0_610 (.A(b[21]), .ZN(n_0_527));
   INV_X1 i_0_611 (.A(b[22]), .ZN(n_0_528));
   INV_X1 i_0_612 (.A(b[23]), .ZN(n_0_529));
   INV_X1 i_0_613 (.A(b[24]), .ZN(n_0_530));
   INV_X1 i_0_614 (.A(b[25]), .ZN(n_0_531));
   INV_X1 i_0_615 (.A(b[26]), .ZN(n_0_532));
   INV_X1 i_0_616 (.A(b[27]), .ZN(n_0_533));
   INV_X1 i_0_617 (.A(b[28]), .ZN(n_0_534));
   INV_X1 i_0_618 (.A(b[29]), .ZN(n_0_535));
   INV_X1 i_0_619 (.A(b[30]), .ZN(n_0_536));
endmodule

module fpa(A, B, O, OF);
   input [31:0]A;
   input [31:0]B;
   output [31:0]O;
   output OF;

   wire OF_adder;
   wire [31:0]adder_out;
   wire [31:0]adder_b_in;
   wire [31:0]adder_a_in;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;

   adder A1 (.a(adder_a_in), .b(adder_b_in), .out(adder_out), .of(OF_adder));
   DLH_X1 \adder_b_in_reg[31]  (.D(B[31]), .G(n_0_0), .Q(adder_b_in[31]));
   DLH_X1 \adder_b_in_reg[30]  (.D(B[30]), .G(n_0_0), .Q(adder_b_in[30]));
   DLH_X1 \adder_b_in_reg[29]  (.D(B[29]), .G(n_0_0), .Q(adder_b_in[29]));
   DLH_X1 \adder_b_in_reg[28]  (.D(B[28]), .G(n_0_0), .Q(adder_b_in[28]));
   DLH_X1 \adder_b_in_reg[27]  (.D(B[27]), .G(n_0_0), .Q(adder_b_in[27]));
   DLH_X1 \adder_b_in_reg[26]  (.D(B[26]), .G(n_0_0), .Q(adder_b_in[26]));
   DLH_X1 \adder_b_in_reg[25]  (.D(B[25]), .G(n_0_0), .Q(adder_b_in[25]));
   DLH_X1 \adder_b_in_reg[24]  (.D(B[24]), .G(n_0_0), .Q(adder_b_in[24]));
   DLH_X1 \adder_b_in_reg[23]  (.D(B[23]), .G(n_0_0), .Q(adder_b_in[23]));
   DLH_X1 \adder_b_in_reg[22]  (.D(B[22]), .G(n_0_0), .Q(adder_b_in[22]));
   DLH_X1 \adder_b_in_reg[21]  (.D(B[21]), .G(n_0_0), .Q(adder_b_in[21]));
   DLH_X1 \adder_b_in_reg[20]  (.D(B[20]), .G(n_0_0), .Q(adder_b_in[20]));
   DLH_X1 \adder_b_in_reg[19]  (.D(B[19]), .G(n_0_0), .Q(adder_b_in[19]));
   DLH_X1 \adder_b_in_reg[18]  (.D(B[18]), .G(n_0_0), .Q(adder_b_in[18]));
   DLH_X1 \adder_b_in_reg[17]  (.D(B[17]), .G(n_0_0), .Q(adder_b_in[17]));
   DLH_X1 \adder_b_in_reg[16]  (.D(B[16]), .G(n_0_0), .Q(adder_b_in[16]));
   DLH_X1 \adder_b_in_reg[15]  (.D(B[15]), .G(n_0_0), .Q(adder_b_in[15]));
   DLH_X1 \adder_b_in_reg[14]  (.D(B[14]), .G(n_0_0), .Q(adder_b_in[14]));
   DLH_X1 \adder_b_in_reg[13]  (.D(B[13]), .G(n_0_0), .Q(adder_b_in[13]));
   DLH_X1 \adder_b_in_reg[12]  (.D(B[12]), .G(n_0_0), .Q(adder_b_in[12]));
   DLH_X1 \adder_b_in_reg[11]  (.D(B[11]), .G(n_0_0), .Q(adder_b_in[11]));
   DLH_X1 \adder_b_in_reg[10]  (.D(B[10]), .G(n_0_0), .Q(adder_b_in[10]));
   DLH_X1 \adder_b_in_reg[9]  (.D(B[9]), .G(n_0_0), .Q(adder_b_in[9]));
   DLH_X1 \adder_b_in_reg[8]  (.D(B[8]), .G(n_0_0), .Q(adder_b_in[8]));
   DLH_X1 \adder_b_in_reg[7]  (.D(B[7]), .G(n_0_0), .Q(adder_b_in[7]));
   DLH_X1 \adder_b_in_reg[6]  (.D(B[6]), .G(n_0_0), .Q(adder_b_in[6]));
   DLH_X1 \adder_b_in_reg[5]  (.D(B[5]), .G(n_0_0), .Q(adder_b_in[5]));
   DLH_X1 \adder_b_in_reg[4]  (.D(B[4]), .G(n_0_0), .Q(adder_b_in[4]));
   DLH_X1 \adder_b_in_reg[3]  (.D(B[3]), .G(n_0_0), .Q(adder_b_in[3]));
   DLH_X1 \adder_b_in_reg[2]  (.D(B[2]), .G(n_0_0), .Q(adder_b_in[2]));
   DLH_X1 \adder_b_in_reg[1]  (.D(B[1]), .G(n_0_0), .Q(adder_b_in[1]));
   DLH_X1 \adder_b_in_reg[0]  (.D(B[0]), .G(n_0_0), .Q(adder_b_in[0]));
   DLH_X1 \adder_a_in_reg[31]  (.D(A[31]), .G(n_0_0), .Q(adder_a_in[31]));
   DLH_X1 \adder_a_in_reg[30]  (.D(A[30]), .G(n_0_0), .Q(adder_a_in[30]));
   DLH_X1 \adder_a_in_reg[29]  (.D(A[29]), .G(n_0_0), .Q(adder_a_in[29]));
   DLH_X1 \adder_a_in_reg[28]  (.D(A[28]), .G(n_0_0), .Q(adder_a_in[28]));
   DLH_X1 \adder_a_in_reg[27]  (.D(A[27]), .G(n_0_0), .Q(adder_a_in[27]));
   DLH_X1 \adder_a_in_reg[26]  (.D(A[26]), .G(n_0_0), .Q(adder_a_in[26]));
   DLH_X1 \adder_a_in_reg[25]  (.D(A[25]), .G(n_0_0), .Q(adder_a_in[25]));
   DLH_X1 \adder_a_in_reg[24]  (.D(A[24]), .G(n_0_0), .Q(adder_a_in[24]));
   DLH_X1 \adder_a_in_reg[23]  (.D(A[23]), .G(n_0_0), .Q(adder_a_in[23]));
   DLH_X1 \adder_a_in_reg[22]  (.D(A[22]), .G(n_0_0), .Q(adder_a_in[22]));
   DLH_X1 \adder_a_in_reg[21]  (.D(A[21]), .G(n_0_0), .Q(adder_a_in[21]));
   DLH_X1 \adder_a_in_reg[20]  (.D(A[20]), .G(n_0_0), .Q(adder_a_in[20]));
   DLH_X1 \adder_a_in_reg[19]  (.D(A[19]), .G(n_0_0), .Q(adder_a_in[19]));
   DLH_X1 \adder_a_in_reg[18]  (.D(A[18]), .G(n_0_0), .Q(adder_a_in[18]));
   DLH_X1 \adder_a_in_reg[17]  (.D(A[17]), .G(n_0_0), .Q(adder_a_in[17]));
   DLH_X1 \adder_a_in_reg[16]  (.D(A[16]), .G(n_0_0), .Q(adder_a_in[16]));
   DLH_X1 \adder_a_in_reg[15]  (.D(A[15]), .G(n_0_0), .Q(adder_a_in[15]));
   DLH_X1 \adder_a_in_reg[14]  (.D(A[14]), .G(n_0_0), .Q(adder_a_in[14]));
   DLH_X1 \adder_a_in_reg[13]  (.D(A[13]), .G(n_0_0), .Q(adder_a_in[13]));
   DLH_X1 \adder_a_in_reg[12]  (.D(A[12]), .G(n_0_0), .Q(adder_a_in[12]));
   DLH_X1 \adder_a_in_reg[11]  (.D(A[11]), .G(n_0_0), .Q(adder_a_in[11]));
   DLH_X1 \adder_a_in_reg[10]  (.D(A[10]), .G(n_0_0), .Q(adder_a_in[10]));
   DLH_X1 \adder_a_in_reg[9]  (.D(A[9]), .G(n_0_0), .Q(adder_a_in[9]));
   DLH_X1 \adder_a_in_reg[8]  (.D(A[8]), .G(n_0_0), .Q(adder_a_in[8]));
   DLH_X1 \adder_a_in_reg[7]  (.D(A[7]), .G(n_0_0), .Q(adder_a_in[7]));
   DLH_X1 \adder_a_in_reg[6]  (.D(A[6]), .G(n_0_0), .Q(adder_a_in[6]));
   DLH_X1 \adder_a_in_reg[5]  (.D(A[5]), .G(n_0_0), .Q(adder_a_in[5]));
   DLH_X1 \adder_a_in_reg[4]  (.D(A[4]), .G(n_0_0), .Q(adder_a_in[4]));
   DLH_X1 \adder_a_in_reg[3]  (.D(A[3]), .G(n_0_0), .Q(adder_a_in[3]));
   DLH_X1 \adder_a_in_reg[2]  (.D(A[2]), .G(n_0_0), .Q(adder_a_in[2]));
   DLH_X1 \adder_a_in_reg[1]  (.D(A[1]), .G(n_0_0), .Q(adder_a_in[1]));
   DLH_X1 \adder_a_in_reg[0]  (.D(A[0]), .G(n_0_0), .Q(adder_a_in[0]));
   AND2_X1 i_0_0_0 (.A1(OF_adder), .A2(n_0_0), .ZN(OF));
   INV_X1 i_0_0_1 (.A(n_0_0_0), .ZN(O[0]));
   AOI222_X1 i_0_0_2 (.A1(adder_out[0]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[0]), 
      .C1(A[0]), .C2(n_0_0_51), .ZN(n_0_0_0));
   INV_X1 i_0_0_3 (.A(n_0_0_1), .ZN(O[1]));
   AOI222_X1 i_0_0_4 (.A1(adder_out[1]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[1]), 
      .C1(A[1]), .C2(n_0_0_51), .ZN(n_0_0_1));
   INV_X1 i_0_0_5 (.A(n_0_0_2), .ZN(O[2]));
   AOI222_X1 i_0_0_6 (.A1(adder_out[2]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[2]), 
      .C1(A[2]), .C2(n_0_0_51), .ZN(n_0_0_2));
   INV_X1 i_0_0_7 (.A(n_0_0_3), .ZN(O[3]));
   AOI222_X1 i_0_0_8 (.A1(adder_out[3]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[3]), 
      .C1(A[3]), .C2(n_0_0_51), .ZN(n_0_0_3));
   INV_X1 i_0_0_9 (.A(n_0_0_4), .ZN(O[4]));
   AOI222_X1 i_0_0_10 (.A1(adder_out[4]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[4]), 
      .C1(A[4]), .C2(n_0_0_51), .ZN(n_0_0_4));
   INV_X1 i_0_0_11 (.A(n_0_0_5), .ZN(O[5]));
   AOI222_X1 i_0_0_12 (.A1(adder_out[5]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[5]), 
      .C1(A[5]), .C2(n_0_0_51), .ZN(n_0_0_5));
   INV_X1 i_0_0_13 (.A(n_0_0_6), .ZN(O[6]));
   AOI222_X1 i_0_0_14 (.A1(adder_out[6]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[6]), 
      .C1(A[6]), .C2(n_0_0_51), .ZN(n_0_0_6));
   INV_X1 i_0_0_15 (.A(n_0_0_7), .ZN(O[7]));
   AOI222_X1 i_0_0_16 (.A1(adder_out[7]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[7]), 
      .C1(A[7]), .C2(n_0_0_51), .ZN(n_0_0_7));
   INV_X1 i_0_0_17 (.A(n_0_0_8), .ZN(O[8]));
   AOI222_X1 i_0_0_18 (.A1(adder_out[8]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[8]), 
      .C1(A[8]), .C2(n_0_0_51), .ZN(n_0_0_8));
   INV_X1 i_0_0_19 (.A(n_0_0_9), .ZN(O[9]));
   AOI222_X1 i_0_0_20 (.A1(adder_out[9]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[9]), 
      .C1(A[9]), .C2(n_0_0_51), .ZN(n_0_0_9));
   INV_X1 i_0_0_21 (.A(n_0_0_10), .ZN(O[10]));
   AOI222_X1 i_0_0_22 (.A1(adder_out[10]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[10]), 
      .C1(A[10]), .C2(n_0_0_51), .ZN(n_0_0_10));
   INV_X1 i_0_0_23 (.A(n_0_0_11), .ZN(O[11]));
   AOI222_X1 i_0_0_24 (.A1(adder_out[11]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[11]), 
      .C1(A[11]), .C2(n_0_0_51), .ZN(n_0_0_11));
   INV_X1 i_0_0_25 (.A(n_0_0_12), .ZN(O[12]));
   AOI222_X1 i_0_0_26 (.A1(adder_out[12]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[12]), 
      .C1(A[12]), .C2(n_0_0_51), .ZN(n_0_0_12));
   INV_X1 i_0_0_27 (.A(n_0_0_13), .ZN(O[13]));
   AOI222_X1 i_0_0_28 (.A1(adder_out[13]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[13]), 
      .C1(A[13]), .C2(n_0_0_51), .ZN(n_0_0_13));
   INV_X1 i_0_0_29 (.A(n_0_0_14), .ZN(O[14]));
   AOI222_X1 i_0_0_30 (.A1(adder_out[14]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[14]), 
      .C1(A[14]), .C2(n_0_0_51), .ZN(n_0_0_14));
   INV_X1 i_0_0_31 (.A(n_0_0_15), .ZN(O[15]));
   AOI222_X1 i_0_0_32 (.A1(adder_out[15]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[15]), 
      .C1(A[15]), .C2(n_0_0_51), .ZN(n_0_0_15));
   INV_X1 i_0_0_33 (.A(n_0_0_16), .ZN(O[16]));
   AOI222_X1 i_0_0_34 (.A1(adder_out[16]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[16]), 
      .C1(A[16]), .C2(n_0_0_51), .ZN(n_0_0_16));
   INV_X1 i_0_0_35 (.A(n_0_0_17), .ZN(O[17]));
   AOI222_X1 i_0_0_36 (.A1(adder_out[17]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[17]), 
      .C1(A[17]), .C2(n_0_0_51), .ZN(n_0_0_17));
   INV_X1 i_0_0_37 (.A(n_0_0_18), .ZN(O[18]));
   AOI222_X1 i_0_0_38 (.A1(adder_out[18]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[18]), 
      .C1(A[18]), .C2(n_0_0_51), .ZN(n_0_0_18));
   INV_X1 i_0_0_39 (.A(n_0_0_19), .ZN(O[19]));
   AOI222_X1 i_0_0_40 (.A1(adder_out[19]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[19]), 
      .C1(A[19]), .C2(n_0_0_51), .ZN(n_0_0_19));
   INV_X1 i_0_0_41 (.A(n_0_0_20), .ZN(O[20]));
   AOI222_X1 i_0_0_42 (.A1(adder_out[20]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[20]), 
      .C1(A[20]), .C2(n_0_0_51), .ZN(n_0_0_20));
   INV_X1 i_0_0_43 (.A(n_0_0_21), .ZN(O[21]));
   AOI222_X1 i_0_0_44 (.A1(adder_out[21]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[21]), 
      .C1(A[21]), .C2(n_0_0_51), .ZN(n_0_0_21));
   INV_X1 i_0_0_45 (.A(n_0_0_22), .ZN(O[22]));
   AOI222_X1 i_0_0_46 (.A1(adder_out[22]), .A2(n_0_0), .B1(n_0_0_32), .B2(B[22]), 
      .C1(A[22]), .C2(n_0_0_51), .ZN(n_0_0_22));
   AOI21_X1 i_0_0_47 (.A(n_0_0_23), .B1(n_0_0_32), .B2(n_0_0_64), .ZN(O[23]));
   OAI22_X1 i_0_0_48 (.A1(n_0_0_33), .A2(adder_out[23]), .B1(A[23]), .B2(
      n_0_0_50), .ZN(n_0_0_23));
   AOI21_X1 i_0_0_49 (.A(n_0_0_24), .B1(n_0_0_32), .B2(n_0_0_65), .ZN(O[24]));
   OAI22_X1 i_0_0_50 (.A1(n_0_0_33), .A2(adder_out[24]), .B1(A[24]), .B2(
      n_0_0_50), .ZN(n_0_0_24));
   AOI21_X1 i_0_0_51 (.A(n_0_0_25), .B1(n_0_0_32), .B2(n_0_0_66), .ZN(O[25]));
   OAI22_X1 i_0_0_52 (.A1(n_0_0_33), .A2(adder_out[25]), .B1(A[25]), .B2(
      n_0_0_50), .ZN(n_0_0_25));
   AOI21_X1 i_0_0_53 (.A(n_0_0_26), .B1(n_0_0_32), .B2(n_0_0_67), .ZN(O[26]));
   OAI22_X1 i_0_0_54 (.A1(n_0_0_33), .A2(adder_out[26]), .B1(A[26]), .B2(
      n_0_0_50), .ZN(n_0_0_26));
   AOI21_X1 i_0_0_55 (.A(n_0_0_27), .B1(n_0_0_32), .B2(n_0_0_68), .ZN(O[27]));
   OAI22_X1 i_0_0_56 (.A1(n_0_0_33), .A2(adder_out[27]), .B1(A[27]), .B2(
      n_0_0_50), .ZN(n_0_0_27));
   AOI21_X1 i_0_0_57 (.A(n_0_0_28), .B1(n_0_0_32), .B2(n_0_0_69), .ZN(O[28]));
   OAI22_X1 i_0_0_58 (.A1(n_0_0_33), .A2(adder_out[28]), .B1(A[28]), .B2(
      n_0_0_50), .ZN(n_0_0_28));
   AOI21_X1 i_0_0_59 (.A(n_0_0_29), .B1(n_0_0_32), .B2(n_0_0_70), .ZN(O[29]));
   OAI22_X1 i_0_0_60 (.A1(n_0_0_33), .A2(adder_out[29]), .B1(A[29]), .B2(
      n_0_0_50), .ZN(n_0_0_29));
   AOI21_X1 i_0_0_61 (.A(n_0_0_30), .B1(n_0_0_32), .B2(n_0_0_71), .ZN(O[30]));
   OAI22_X1 i_0_0_62 (.A1(n_0_0_33), .A2(adder_out[30]), .B1(A[30]), .B2(
      n_0_0_50), .ZN(n_0_0_30));
   AOI21_X1 i_0_0_63 (.A(n_0_0_31), .B1(n_0_0_32), .B2(n_0_0_72), .ZN(O[31]));
   OAI22_X1 i_0_0_64 (.A1(n_0_0_33), .A2(adder_out[31]), .B1(A[31]), .B2(
      n_0_0_50), .ZN(n_0_0_31));
   NOR2_X1 i_0_0_65 (.A1(n_0_0_34), .A2(n_0_0_51), .ZN(n_0_0_32));
   INV_X1 i_0_0_66 (.A(n_0_0_33), .ZN(n_0_0));
   NAND2_X1 i_0_0_67 (.A1(n_0_0_50), .A2(n_0_0_34), .ZN(n_0_0_33));
   NOR2_X1 i_0_0_68 (.A1(n_0_0_38), .A2(n_0_0_35), .ZN(n_0_0_34));
   NOR2_X1 i_0_0_69 (.A1(n_0_0_37), .A2(n_0_0_36), .ZN(n_0_0_35));
   NAND4_X1 i_0_0_70 (.A1(B[30]), .A2(B[29]), .A3(B[28]), .A4(B[27]), .ZN(
      n_0_0_36));
   NAND4_X1 i_0_0_71 (.A1(B[26]), .A2(B[25]), .A3(B[24]), .A4(B[23]), .ZN(
      n_0_0_37));
   NOR4_X1 i_0_0_72 (.A1(n_0_0_46), .A2(n_0_0_44), .A3(n_0_0_41), .A4(n_0_0_39), 
      .ZN(n_0_0_38));
   NAND3_X1 i_0_0_73 (.A1(n_0_0_45), .A2(n_0_0_43), .A3(n_0_0_40), .ZN(n_0_0_39));
   NOR4_X1 i_0_0_74 (.A1(n_0_0_47), .A2(A[1]), .A3(A[4]), .A4(A[5]), .ZN(
      n_0_0_40));
   NAND3_X1 i_0_0_75 (.A1(n_0_0_49), .A2(n_0_0_48), .A3(n_0_0_42), .ZN(n_0_0_41));
   NOR4_X1 i_0_0_76 (.A1(A[6]), .A2(A[3]), .A3(A[2]), .A4(A[0]), .ZN(n_0_0_42));
   NOR4_X1 i_0_0_77 (.A1(A[18]), .A2(A[17]), .A3(A[16]), .A4(A[15]), .ZN(
      n_0_0_43));
   OR4_X1 i_0_0_78 (.A1(A[22]), .A2(A[21]), .A3(A[20]), .A4(A[19]), .ZN(n_0_0_44));
   NOR4_X1 i_0_0_79 (.A1(A[30]), .A2(A[29]), .A3(A[28]), .A4(A[27]), .ZN(
      n_0_0_45));
   OR4_X1 i_0_0_80 (.A1(A[26]), .A2(A[25]), .A3(A[24]), .A4(A[23]), .ZN(n_0_0_46));
   OR4_X1 i_0_0_81 (.A1(A[14]), .A2(A[13]), .A3(A[12]), .A4(A[11]), .ZN(n_0_0_47));
   NOR2_X1 i_0_0_82 (.A1(A[10]), .A2(A[7]), .ZN(n_0_0_48));
   NOR2_X1 i_0_0_83 (.A1(A[9]), .A2(A[8]), .ZN(n_0_0_49));
   INV_X1 i_0_0_84 (.A(n_0_0_51), .ZN(n_0_0_50));
   OAI22_X1 i_0_0_85 (.A1(n_0_0_56), .A2(n_0_0_54), .B1(n_0_0_53), .B2(n_0_0_52), 
      .ZN(n_0_0_51));
   NAND4_X1 i_0_0_86 (.A1(A[30]), .A2(A[29]), .A3(A[28]), .A4(A[27]), .ZN(
      n_0_0_52));
   NAND4_X1 i_0_0_87 (.A1(A[26]), .A2(A[25]), .A3(A[24]), .A4(A[23]), .ZN(
      n_0_0_53));
   NAND3_X1 i_0_0_88 (.A1(n_0_0_60), .A2(n_0_0_58), .A3(n_0_0_55), .ZN(n_0_0_54));
   NOR4_X1 i_0_0_89 (.A1(n_0_0_62), .A2(B[1]), .A3(B[4]), .A4(B[5]), .ZN(
      n_0_0_55));
   NAND4_X1 i_0_0_90 (.A1(n_0_0_63), .A2(n_0_0_61), .A3(n_0_0_59), .A4(n_0_0_57), 
      .ZN(n_0_0_56));
   NOR4_X1 i_0_0_91 (.A1(B[6]), .A2(B[3]), .A3(B[2]), .A4(B[0]), .ZN(n_0_0_57));
   NOR4_X1 i_0_0_92 (.A1(B[18]), .A2(B[17]), .A3(B[16]), .A4(B[15]), .ZN(
      n_0_0_58));
   NOR4_X1 i_0_0_93 (.A1(B[22]), .A2(B[21]), .A3(B[20]), .A4(B[19]), .ZN(
      n_0_0_59));
   NOR4_X1 i_0_0_94 (.A1(B[30]), .A2(B[29]), .A3(B[28]), .A4(B[27]), .ZN(
      n_0_0_60));
   NOR4_X1 i_0_0_95 (.A1(B[26]), .A2(B[25]), .A3(B[24]), .A4(B[23]), .ZN(
      n_0_0_61));
   OR4_X1 i_0_0_96 (.A1(B[14]), .A2(B[13]), .A3(B[12]), .A4(B[11]), .ZN(n_0_0_62));
   NOR4_X1 i_0_0_97 (.A1(B[10]), .A2(B[9]), .A3(B[8]), .A4(B[7]), .ZN(n_0_0_63));
   INV_X1 i_0_0_98 (.A(B[23]), .ZN(n_0_0_64));
   INV_X1 i_0_0_99 (.A(B[24]), .ZN(n_0_0_65));
   INV_X1 i_0_0_100 (.A(B[25]), .ZN(n_0_0_66));
   INV_X1 i_0_0_101 (.A(B[26]), .ZN(n_0_0_67));
   INV_X1 i_0_0_102 (.A(B[27]), .ZN(n_0_0_68));
   INV_X1 i_0_0_103 (.A(B[28]), .ZN(n_0_0_69));
   INV_X1 i_0_0_104 (.A(B[29]), .ZN(n_0_0_70));
   INV_X1 i_0_0_105 (.A(B[30]), .ZN(n_0_0_71));
   INV_X1 i_0_0_106 (.A(B[31]), .ZN(n_0_0_72));
endmodule
