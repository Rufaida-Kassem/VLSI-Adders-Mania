/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Nov  4 15:53:13 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1999776946 */

module FullAdder__1_3(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_7(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_11(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_15(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_19(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_23(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_27(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_31(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_35(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_39(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_43(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_47(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_51(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_55(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_59(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_63(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_67(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_71(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_75(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_79(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_83(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_87(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_91(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_95(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_99(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(B), .A2(A), .ZN(Cout));
endmodule

module FullAdder__1_103(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_107(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_111(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_115(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_119(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_123(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_127(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_131(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_135(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_139(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_143(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_147(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_151(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_155(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_159(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_163(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_167(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_171(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_175(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_179(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_183(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder__1_187(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   wire S0;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S0));
   XOR2_X1 i_0_1 (.A(S0), .B(Cin), .Z(S));
   AOI22_X1 i_0_2 (.A1(S0), .A2(Cin), .B1(A), .B2(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(Cout));
endmodule

module FullAdder(A, B, Cin, S, Cout);
   input A;
   input B;
   input Cin;
   output S;
   output Cout;

   XOR2_X1 i_0_0 (.A(B), .B(Cin), .Z(S));
endmodule

module CSA(X, Y, Cin, S, Cout, OF);
   input [23:0]X;
   input [23:0]Y;
   input Cin;
   output [23:0]S;
   output Cout;
   output OF;

   wire Cout0;
   wire Cin1;

   FullAdder__1_3 genblk1_0_FA (.A(X[0]), .B(Y[0]), .Cin(), .S(S[0]), .Cout(
      Cout0));
   FullAdder__1_7 genblk1_1_FA (.A(X[1]), .B(Y[1]), .Cin(), .S(n_1), .Cout(n_0));
   FullAdder__1_11 genblk1_2_FA (.A(X[2]), .B(Y[2]), .Cin(), .S(n_3), .Cout(n_2));
   FullAdder__1_15 genblk1_3_FA (.A(X[3]), .B(Y[3]), .Cin(), .S(n_5), .Cout(n_4));
   FullAdder__1_19 genblk1_4_FA (.A(X[4]), .B(Y[4]), .Cin(), .S(n_7), .Cout(n_6));
   FullAdder__1_23 genblk1_5_FA (.A(X[5]), .B(Y[5]), .Cin(), .S(n_9), .Cout(n_8));
   FullAdder__1_27 genblk1_6_FA (.A(X[6]), .B(Y[6]), .Cin(), .S(n_11), .Cout(
      n_10));
   FullAdder__1_31 genblk1_7_FA (.A(X[7]), .B(Y[7]), .Cin(), .S(n_13), .Cout(
      n_12));
   FullAdder__1_35 genblk1_8_FA (.A(X[8]), .B(Y[8]), .Cin(), .S(n_15), .Cout(
      n_14));
   FullAdder__1_39 genblk1_9_FA (.A(X[9]), .B(Y[9]), .Cin(), .S(n_17), .Cout(
      n_16));
   FullAdder__1_43 genblk1_10_FA (.A(X[10]), .B(Y[10]), .Cin(), .S(n_19), 
      .Cout(n_18));
   FullAdder__1_47 genblk1_11_FA (.A(X[11]), .B(Y[11]), .Cin(), .S(n_21), 
      .Cout(n_20));
   FullAdder__1_51 genblk1_12_FA (.A(X[12]), .B(Y[12]), .Cin(), .S(n_23), 
      .Cout(n_22));
   FullAdder__1_55 genblk1_13_FA (.A(X[13]), .B(Y[13]), .Cin(), .S(n_25), 
      .Cout(n_24));
   FullAdder__1_59 genblk1_14_FA (.A(X[14]), .B(Y[14]), .Cin(), .S(n_27), 
      .Cout(n_26));
   FullAdder__1_63 genblk1_15_FA (.A(X[15]), .B(Y[15]), .Cin(), .S(n_29), 
      .Cout(n_28));
   FullAdder__1_67 genblk1_16_FA (.A(X[16]), .B(Y[16]), .Cin(), .S(n_31), 
      .Cout(n_30));
   FullAdder__1_71 genblk1_17_FA (.A(X[17]), .B(Y[17]), .Cin(), .S(n_33), 
      .Cout(n_32));
   FullAdder__1_75 genblk1_18_FA (.A(X[18]), .B(Y[18]), .Cin(), .S(n_35), 
      .Cout(n_34));
   FullAdder__1_79 genblk1_19_FA (.A(X[19]), .B(Y[19]), .Cin(), .S(n_37), 
      .Cout(n_36));
   FullAdder__1_83 genblk1_20_FA (.A(X[20]), .B(Y[20]), .Cin(), .S(n_39), 
      .Cout(n_38));
   FullAdder__1_87 genblk1_21_FA (.A(X[21]), .B(Y[21]), .Cin(), .S(n_41), 
      .Cout(n_40));
   FullAdder__1_91 genblk1_22_FA (.A(X[22]), .B(Y[22]), .Cin(), .S(n_43), 
      .Cout(n_42));
   FullAdder__1_95 genblk1_23_FA (.A(X[23]), .B(Y[23]), .Cin(), .S(n_45), 
      .Cout(n_44));
   FullAdder__1_99 genblk2_0_FA (.A(n_1), .B(Cout0), .Cin(), .S(S[1]), .Cout(
      Cin1));
   FullAdder__1_103 genblk2_1_FA (.A(n_3), .B(n_0), .Cin(Cin1), .S(S[2]), 
      .Cout(n_46));
   FullAdder__1_107 genblk2_2_FA (.A(n_5), .B(n_2), .Cin(n_46), .S(S[3]), 
      .Cout(n_47));
   FullAdder__1_111 genblk2_3_FA (.A(n_7), .B(n_4), .Cin(n_47), .S(S[4]), 
      .Cout(n_48));
   FullAdder__1_115 genblk2_4_FA (.A(n_9), .B(n_6), .Cin(n_48), .S(S[5]), 
      .Cout(n_49));
   FullAdder__1_119 genblk2_5_FA (.A(n_11), .B(n_8), .Cin(n_49), .S(S[6]), 
      .Cout(n_50));
   FullAdder__1_123 genblk2_6_FA (.A(n_13), .B(n_10), .Cin(n_50), .S(S[7]), 
      .Cout(n_51));
   FullAdder__1_127 genblk2_7_FA (.A(n_15), .B(n_12), .Cin(n_51), .S(S[8]), 
      .Cout(n_52));
   FullAdder__1_131 genblk2_8_FA (.A(n_17), .B(n_14), .Cin(n_52), .S(S[9]), 
      .Cout(n_53));
   FullAdder__1_135 genblk2_9_FA (.A(n_19), .B(n_16), .Cin(n_53), .S(S[10]), 
      .Cout(n_54));
   FullAdder__1_139 genblk2_10_FA (.A(n_21), .B(n_18), .Cin(n_54), .S(S[11]), 
      .Cout(n_55));
   FullAdder__1_143 genblk2_11_FA (.A(n_23), .B(n_20), .Cin(n_55), .S(S[12]), 
      .Cout(n_56));
   FullAdder__1_147 genblk2_12_FA (.A(n_25), .B(n_22), .Cin(n_56), .S(S[13]), 
      .Cout(n_57));
   FullAdder__1_151 genblk2_13_FA (.A(n_27), .B(n_24), .Cin(n_57), .S(S[14]), 
      .Cout(n_58));
   FullAdder__1_155 genblk2_14_FA (.A(n_29), .B(n_26), .Cin(n_58), .S(S[15]), 
      .Cout(n_59));
   FullAdder__1_159 genblk2_15_FA (.A(n_31), .B(n_28), .Cin(n_59), .S(S[16]), 
      .Cout(n_60));
   FullAdder__1_163 genblk2_16_FA (.A(n_33), .B(n_30), .Cin(n_60), .S(S[17]), 
      .Cout(n_61));
   FullAdder__1_167 genblk2_17_FA (.A(n_35), .B(n_32), .Cin(n_61), .S(S[18]), 
      .Cout(n_62));
   FullAdder__1_171 genblk2_18_FA (.A(n_37), .B(n_34), .Cin(n_62), .S(S[19]), 
      .Cout(n_63));
   FullAdder__1_175 genblk2_19_FA (.A(n_39), .B(n_36), .Cin(n_63), .S(S[20]), 
      .Cout(n_64));
   FullAdder__1_179 genblk2_20_FA (.A(n_41), .B(n_38), .Cin(n_64), .S(S[21]), 
      .Cout(n_65));
   FullAdder__1_183 genblk2_21_FA (.A(n_43), .B(n_40), .Cin(n_65), .S(S[22]), 
      .Cout(n_66));
   FullAdder__1_187 genblk2_22_FA (.A(n_45), .B(n_42), .Cin(n_66), .S(S[23]), 
      .Cout(n_67));
   FullAdder genblk2_23_FA (.A(), .B(n_44), .Cin(n_67), .S(Cout), .Cout());
endmodule

module addition_normaliser(in_e, in_m, out_e, out_m);
   input [7:0]in_e;
   input [24:0]in_m;
   output [7:0]out_e;
   output [24:0]out_m;

   wire n_0_23;
   wire n_0_2;
   wire n_0_24;
   wire n_0_1;
   wire n_0_25;
   wire n_0_0;
   wire n_0_26;
   wire n_0_3;
   wire n_0_27;
   wire n_0_4;
   wire n_0_28;
   wire n_0_5;
   wire n_0_29;
   wire n_0_6;
   wire n_0_30;
   wire n_0_7;
   wire n_0_31;
   wire n_0_8;
   wire n_0_32;
   wire n_0_9;
   wire n_0_33;
   wire n_0_10;
   wire n_0_34;
   wire n_0_11;
   wire n_0_35;
   wire n_0_12;
   wire n_0_36;
   wire n_0_13;
   wire n_0_37;
   wire n_0_14;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_15;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_16;
   wire n_0_17;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_18;
   wire n_0_19;
   wire n_0_167;
   wire n_0_20;
   wire n_0_168;
   wire n_0_21;
   wire n_0_169;
   wire n_0_22;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_317;
   wire n_0_318;
   wire n_0_319;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_332;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_337;
   wire n_0_338;
   wire n_0_339;
   wire n_0_340;
   wire n_0_341;
   wire n_0_342;
   wire n_0_343;
   wire n_0_344;
   wire n_0_345;
   wire n_0_346;
   wire n_0_347;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_355;
   wire n_0_356;
   wire n_0_357;
   wire n_0_358;
   wire n_0_359;
   wire n_0_360;
   wire n_0_361;
   wire n_0_362;
   wire n_0_363;
   wire n_0_364;
   wire n_0_365;
   wire n_0_366;
   wire n_0_367;
   wire n_0_368;
   wire n_0_369;
   wire n_0_370;
   wire n_0_371;
   wire n_0_372;
   wire n_0_373;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_377;
   wire n_0_378;
   wire n_0_379;
   wire n_0_380;
   wire n_0_381;
   wire n_0_382;
   wire n_0_383;
   wire n_0_384;
   wire n_0_385;
   wire n_0_386;
   wire n_0_387;
   wire n_0_388;
   wire n_0_389;
   wire n_0_390;
   wire n_0_391;
   wire n_0_392;
   wire n_0_393;
   wire n_0_394;
   wire n_0_395;
   wire n_0_396;
   wire n_0_397;
   wire n_0_398;
   wire n_0_399;
   wire n_0_400;
   wire n_0_401;
   wire n_0_402;
   wire n_0_403;
   wire n_0_404;
   wire n_0_405;
   wire n_0_406;
   wire n_0_407;
   wire n_0_408;
   wire n_0_409;
   wire n_0_410;
   wire n_0_411;
   wire n_0_412;
   wire n_0_413;
   wire n_0_414;
   wire n_0_415;
   wire n_0_416;
   wire n_0_417;
   wire n_0_418;
   wire n_0_419;
   wire n_0_420;
   wire n_0_421;
   wire n_0_422;
   wire n_0_423;
   wire n_0_424;
   wire n_0_425;
   wire n_0_426;
   wire n_0_427;
   wire n_0_428;
   wire n_0_429;
   wire n_0_430;
   wire n_0_431;
   wire n_0_432;
   wire n_0_433;
   wire n_0_434;
   wire n_0_435;
   wire n_0_436;
   wire n_0_437;
   wire n_0_438;
   wire n_0_439;
   wire n_0_440;
   wire n_0_441;
   wire n_0_442;
   wire n_0_443;
   wire n_0_444;
   wire n_0_445;
   wire n_0_446;
   wire n_0_447;
   wire n_0_448;
   wire n_0_449;
   wire n_0_450;
   wire n_0_451;
   wire n_0_452;
   wire n_0_453;
   wire n_0_454;
   wire n_0_455;
   wire n_0_456;
   wire n_0_457;
   wire n_0_458;
   wire n_0_459;
   wire n_0_460;
   wire n_0_461;
   wire n_0_462;
   wire n_0_463;
   wire n_0_464;
   wire n_0_465;
   wire n_0_466;
   wire n_0_467;
   wire n_0_468;
   wire n_0_469;
   wire n_0_470;
   wire n_0_471;
   wire n_0_472;
   wire n_0_473;
   wire n_0_474;
   wire n_0_475;
   wire n_0_476;
   wire n_0_477;
   wire n_0_478;
   wire n_0_479;
   wire n_0_480;
   wire n_0_481;
   wire n_0_482;
   wire n_0_483;
   wire n_0_484;
   wire n_0_485;
   wire n_0_486;
   wire n_0_487;
   wire n_0_488;
   wire n_0_489;
   wire n_0_490;
   wire n_0_491;
   wire n_0_492;
   wire n_0_493;
   wire n_0_494;
   wire n_0_495;
   wire n_0_496;
   wire n_0_497;
   wire n_0_498;
   wire n_0_499;
   wire n_0_500;
   wire n_0_501;
   wire n_0_502;
   wire n_0_503;
   wire n_0_504;
   wire n_0_505;
   wire n_0_506;
   wire n_0_507;
   wire n_0_508;
   wire n_0_509;
   wire n_0_510;
   wire n_0_511;
   wire n_0_512;
   wire n_0_513;
   wire n_0_514;
   wire n_0_515;
   wire n_0_516;
   wire n_0_517;

   DLH_X1 \out_m_reg[22]  (.D(n_30), .G(n_8), .Q(out_m[22]));
   DLH_X1 \out_m_reg[21]  (.D(n_29), .G(n_8), .Q(out_m[21]));
   DLH_X1 \out_m_reg[20]  (.D(n_28), .G(n_8), .Q(out_m[20]));
   DLH_X1 \out_m_reg[19]  (.D(n_27), .G(n_8), .Q(out_m[19]));
   DLH_X1 \out_m_reg[18]  (.D(n_26), .G(n_8), .Q(out_m[18]));
   DLH_X1 \out_m_reg[17]  (.D(n_25), .G(n_8), .Q(out_m[17]));
   DLH_X1 \out_m_reg[16]  (.D(n_24), .G(n_8), .Q(out_m[16]));
   DLH_X1 \out_m_reg[15]  (.D(n_23), .G(n_8), .Q(out_m[15]));
   DLH_X1 \out_m_reg[14]  (.D(n_22), .G(n_8), .Q(out_m[14]));
   DLH_X1 \out_m_reg[13]  (.D(n_21), .G(n_8), .Q(out_m[13]));
   DLH_X1 \out_m_reg[12]  (.D(n_20), .G(n_8), .Q(out_m[12]));
   DLH_X1 \out_m_reg[11]  (.D(n_19), .G(n_8), .Q(out_m[11]));
   DLH_X1 \out_m_reg[10]  (.D(n_18), .G(n_8), .Q(out_m[10]));
   DLH_X1 \out_m_reg[9]  (.D(n_17), .G(n_8), .Q(out_m[9]));
   DLH_X1 \out_m_reg[8]  (.D(n_16), .G(n_8), .Q(out_m[8]));
   DLH_X1 \out_m_reg[7]  (.D(n_15), .G(n_8), .Q(out_m[7]));
   DLH_X1 \out_m_reg[6]  (.D(n_14), .G(n_8), .Q(out_m[6]));
   DLH_X1 \out_m_reg[5]  (.D(n_13), .G(n_8), .Q(out_m[5]));
   DLH_X1 \out_m_reg[4]  (.D(n_12), .G(n_8), .Q(out_m[4]));
   DLH_X1 \out_m_reg[3]  (.D(n_11), .G(n_8), .Q(out_m[3]));
   DLH_X1 \out_m_reg[2]  (.D(n_10), .G(n_8), .Q(out_m[2]));
   DLH_X1 \out_m_reg[1]  (.D(n_9), .G(n_8), .Q(out_m[1]));
   DLH_X1 \out_e_reg[7]  (.D(n_7), .G(n_8), .Q(out_e[7]));
   DLH_X1 \out_e_reg[6]  (.D(n_6), .G(n_8), .Q(out_e[6]));
   DLH_X1 \out_e_reg[5]  (.D(n_5), .G(n_8), .Q(out_e[5]));
   DLH_X1 \out_e_reg[4]  (.D(n_4), .G(n_8), .Q(out_e[4]));
   DLH_X1 \out_e_reg[3]  (.D(n_3), .G(n_8), .Q(out_e[3]));
   DLH_X1 \out_e_reg[2]  (.D(n_2), .G(n_8), .Q(out_e[2]));
   DLH_X1 \out_e_reg[1]  (.D(n_1), .G(n_8), .Q(out_e[1]));
   DLH_X1 \out_e_reg[0]  (.D(n_0), .G(n_8), .Q(out_e[0]));
   HA_X1 i_0_0 (.A(in_e[3]), .B(n_0_15), .CO(n_0_2), .S(n_0_23));
   HA_X1 i_0_1 (.A(in_e[3]), .B(n_0_19), .CO(n_0_1), .S(n_0_24));
   HA_X1 i_0_2 (.A(in_e[3]), .B(n_0_22), .CO(n_0_0), .S(n_0_25));
   HA_X1 i_0_3 (.A(in_e[3]), .B(in_e[2]), .CO(n_0_3), .S(n_0_26));
   HA_X1 i_0_4 (.A(in_e[3]), .B(n_0_12), .CO(n_0_4), .S(n_0_27));
   HA_X1 i_0_5 (.A(in_e[3]), .B(n_0_13), .CO(n_0_5), .S(n_0_28));
   HA_X1 i_0_6 (.A(in_e[3]), .B(n_0_14), .CO(n_0_6), .S(n_0_29));
   HA_X1 i_0_7 (.A(in_e[4]), .B(n_0_16), .CO(n_0_7), .S(n_0_30));
   HA_X1 i_0_8 (.A(in_e[4]), .B(n_0_18), .CO(n_0_8), .S(n_0_31));
   HA_X1 i_0_9 (.A(in_e[4]), .B(n_0_20), .CO(n_0_9), .S(n_0_32));
   HA_X1 i_0_10 (.A(in_e[4]), .B(n_0_21), .CO(n_0_10), .S(n_0_33));
   HA_X1 i_0_11 (.A(in_e[1]), .B(in_e[0]), .CO(n_0_11), .S(n_0_34));
   HA_X1 i_0_12 (.A(in_e[2]), .B(n_0_17), .CO(n_0_12), .S(n_0_35));
   HA_X1 i_0_13 (.A(in_e[2]), .B(in_e[1]), .CO(n_0_13), .S(n_0_36));
   HA_X1 i_0_14 (.A(in_e[2]), .B(n_0_11), .CO(n_0_14), .S(n_0_37));
   XOR2_X1 i_0_15 (.A(in_e[0]), .B(n_0_38), .Z(n_0));
   AOI211_X1 i_0_16 (.A(n_0_403), .B(n_0_39), .C1(n_0_181), .C2(n_0_41), 
      .ZN(n_0_38));
   AOI211_X1 i_0_17 (.A(n_0_480), .B(n_0_375), .C1(n_0_509), .C2(n_0_40), 
      .ZN(n_0_39));
   OAI22_X1 i_0_18 (.A1(in_m[19]), .A2(n_0_508), .B1(n_0_393), .B2(n_0_192), 
      .ZN(n_0_40));
   NAND3_X1 i_0_19 (.A1(n_0_503), .A2(n_0_312), .A3(n_0_42), .ZN(n_0_41));
   OAI211_X1 i_0_20 (.A(n_0_502), .B(n_0_500), .C1(n_0_151), .C2(n_0_59), 
      .ZN(n_0_42));
   OAI221_X1 i_0_21 (.A(n_0_43), .B1(n_0_514), .B2(n_0_54), .C1(n_0_66), 
      .C2(n_0_63), .ZN(n_1));
   AOI221_X1 i_0_22 (.A(n_0_49), .B1(n_0_514), .B2(n_0_403), .C1(n_0_34), 
      .C2(n_0_44), .ZN(n_0_43));
   OAI21_X1 i_0_23 (.A(n_0_45), .B1(n_0_172), .B2(n_0_46), .ZN(n_0_44));
   AOI21_X1 i_0_24 (.A(n_0_464), .B1(n_0_510), .B2(n_0_47), .ZN(n_0_45));
   AOI21_X1 i_0_25 (.A(n_0_53), .B1(in_e[1]), .B2(n_0_194), .ZN(n_0_46));
   AOI21_X1 i_0_26 (.A(n_0_508), .B1(n_0_65), .B2(n_0_48), .ZN(n_0_47));
   NAND3_X1 i_0_27 (.A1(in_e[1]), .A2(n_0_471), .A3(n_0_509), .ZN(n_0_48));
   AOI21_X1 i_0_28 (.A(n_0_109), .B1(n_0_484), .B2(n_0_50), .ZN(n_0_49));
   INV_X1 i_0_29 (.A(n_0_51), .ZN(n_0_50));
   OAI33_X1 i_0_30 (.A1(n_0_514), .A2(n_0_195), .A3(n_0_197), .B1(n_0_186), 
      .B2(n_0_52), .B3(n_0_380), .ZN(n_0_51));
   NAND3_X1 i_0_31 (.A1(n_0_510), .A2(n_0_508), .A3(n_0_53), .ZN(n_0_52));
   NOR2_X1 i_0_32 (.A1(in_e[1]), .A2(n_0_192), .ZN(n_0_53));
   AOI21_X1 i_0_33 (.A(n_0_55), .B1(n_0_477), .B2(n_0_60), .ZN(n_0_54));
   AOI211_X1 i_0_34 (.A(n_0_195), .B(n_0_182), .C1(n_0_57), .C2(n_0_56), 
      .ZN(n_0_55));
   AOI221_X1 i_0_35 (.A(in_m[11]), .B1(in_m[10]), .B2(n_0_108), .C1(n_0_343), 
      .C2(n_0_58), .ZN(n_0_56));
   OAI211_X1 i_0_36 (.A(n_0_34), .B(n_0_437), .C1(in_m[8]), .C2(n_0_357), 
      .ZN(n_0_57));
   OAI211_X1 i_0_37 (.A(n_0_499), .B(n_0_130), .C1(n_0_498), .C2(n_0_109), 
      .ZN(n_0_58));
   NAND2_X1 i_0_38 (.A1(n_0_499), .A2(n_0_130), .ZN(n_0_59));
   OAI221_X1 i_0_39 (.A(n_0_511), .B1(n_0_510), .B2(n_0_109), .C1(n_0_62), 
      .C2(n_0_61), .ZN(n_0_60));
   NAND2_X1 i_0_40 (.A1(n_0_509), .A2(n_0_508), .ZN(n_0_61));
   AOI22_X1 i_0_41 (.A1(in_m[14]), .A2(n_0_108), .B1(n_0_510), .B2(in_m[15]), 
      .ZN(n_0_62));
   INV_X1 i_0_42 (.A(n_0_64), .ZN(n_0_63));
   AOI21_X1 i_0_43 (.A(n_0_65), .B1(in_e[0]), .B2(in_m[18]), .ZN(n_0_64));
   NAND3_X1 i_0_44 (.A1(n_0_514), .A2(n_0_511), .A3(n_0_479), .ZN(n_0_65));
   NOR3_X1 i_0_45 (.A1(in_m[18]), .A2(in_m[17]), .A3(n_0_67), .ZN(n_0_66));
   AOI211_X1 i_0_46 (.A(in_m[16]), .B(in_m[15]), .C1(n_0_70), .C2(n_0_68), 
      .ZN(n_0_67));
   AOI211_X1 i_0_47 (.A(n_0_393), .B(n_0_69), .C1(in_m[14]), .C2(n_0_108), 
      .ZN(n_0_68));
   AND3_X1 i_0_48 (.A1(in_m[10]), .A2(n_0_108), .A3(n_0_434), .ZN(n_0_69));
   NAND3_X1 i_0_49 (.A1(n_0_502), .A2(n_0_379), .A3(n_0_71), .ZN(n_0_70));
   NAND2_X1 i_0_50 (.A1(n_0_501), .A2(n_0_72), .ZN(n_0_71));
   AOI22_X1 i_0_51 (.A1(in_m[8]), .A2(n_0_34), .B1(n_0_499), .B2(n_0_73), 
      .ZN(n_0_72));
   AOI21_X1 i_0_52 (.A(n_0_74), .B1(in_m[6]), .B2(n_0_109), .ZN(n_0_73));
   AOI22_X1 i_0_53 (.A1(n_0_500), .A2(n_0_360), .B1(in_m[4]), .B2(n_0_34), 
      .ZN(n_0_74));
   NAND4_X1 i_0_54 (.A1(n_0_85), .A2(n_0_83), .A3(n_0_80), .A4(n_0_75), .ZN(n_2));
   AOI22_X1 i_0_55 (.A1(n_0_91), .A2(n_0_90), .B1(n_0_77), .B2(n_0_76), .ZN(
      n_0_75));
   OAI21_X1 i_0_56 (.A(n_0_15), .B1(n_0_515), .B2(n_0_157), .ZN(n_0_76));
   INV_X1 i_0_57 (.A(n_0_78), .ZN(n_0_77));
   AOI21_X1 i_0_58 (.A(n_0_483), .B1(n_0_196), .B2(n_0_79), .ZN(n_0_78));
   OAI22_X1 i_0_59 (.A1(in_m[7]), .A2(n_0_100), .B1(in_m[3]), .B2(n_0_98), 
      .ZN(n_0_79));
   AOI22_X1 i_0_60 (.A1(in_e[2]), .A2(n_0_86), .B1(n_0_515), .B2(n_0_81), 
      .ZN(n_0_80));
   OAI221_X1 i_0_61 (.A(n_0_402), .B1(in_e[1]), .B2(n_0_404), .C1(n_0_451), 
      .C2(n_0_82), .ZN(n_0_81));
   NAND2_X1 i_0_62 (.A1(n_0_447), .A2(n_0_89), .ZN(n_0_82));
   AOI222_X1 i_0_63 (.A1(n_0_37), .A2(n_0_308), .B1(n_0_183), .B2(n_0_84), 
      .C1(n_0_464), .C2(n_0_169), .ZN(n_0_83));
   AOI211_X1 i_0_64 (.A(n_0_100), .B(n_0_434), .C1(in_m[12]), .C2(n_0_11), 
      .ZN(n_0_84));
   AOI22_X1 i_0_65 (.A1(n_0_36), .A2(n_0_294), .B1(n_0_35), .B2(n_0_373), 
      .ZN(n_0_85));
   OAI221_X1 i_0_66 (.A(n_0_87), .B1(n_0_514), .B2(n_0_404), .C1(n_0_485), 
      .C2(n_0_465), .ZN(n_0_86));
   OAI21_X1 i_0_67 (.A(n_0_396), .B1(in_m[15]), .B2(n_0_88), .ZN(n_0_87));
   OAI22_X1 i_0_68 (.A1(n_0_368), .A2(n_0_99), .B1(n_0_446), .B2(n_0_89), 
      .ZN(n_0_88));
   AOI21_X1 i_0_69 (.A(in_e[1]), .B1(in_e[0]), .B2(in_m[14]), .ZN(n_0_89));
   AOI21_X1 i_0_70 (.A(n_0_182), .B1(n_0_100), .B2(n_0_98), .ZN(n_0_90));
   OAI221_X1 i_0_71 (.A(n_0_93), .B1(in_m[10]), .B2(n_0_92), .C1(n_0_95), 
      .C2(n_0_94), .ZN(n_0_91));
   AOI22_X1 i_0_72 (.A1(in_m[9]), .A2(n_0_36), .B1(n_0_37), .B2(n_0_281), 
      .ZN(n_0_92));
   NAND2_X1 i_0_73 (.A1(in_m[10]), .A2(n_0_35), .ZN(n_0_93));
   OAI21_X1 i_0_74 (.A(n_0_343), .B1(n_0_499), .B2(n_0_97), .ZN(n_0_94));
   AOI21_X1 i_0_75 (.A(n_0_96), .B1(n_0_360), .B2(n_0_101), .ZN(n_0_95));
   OAI221_X1 i_0_76 (.A(n_0_499), .B1(n_0_130), .B2(n_0_100), .C1(n_0_358), 
      .C2(n_0_99), .ZN(n_0_96));
   INV_X1 i_0_77 (.A(n_0_98), .ZN(n_0_97));
   NAND2_X1 i_0_78 (.A1(in_e[2]), .A2(n_0_193), .ZN(n_0_98));
   AOI21_X1 i_0_79 (.A(n_0_169), .B1(in_e[2]), .B2(n_0_11), .ZN(n_0_99));
   NAND3_X1 i_0_80 (.A1(n_0_515), .A2(n_0_507), .A3(n_0_194), .ZN(n_0_100));
   OAI21_X1 i_0_81 (.A(n_0_106), .B1(n_0_515), .B2(n_0_107), .ZN(n_0_101));
   NAND4_X1 i_0_82 (.A1(n_0_125), .A2(n_0_116), .A3(n_0_113), .A4(n_0_102), 
      .ZN(n_3));
   NAND3_X1 i_0_83 (.A1(n_0_181), .A2(n_0_119), .A3(n_0_103), .ZN(n_0_102));
   INV_X1 i_0_84 (.A(n_0_104), .ZN(n_0_103));
   AOI22_X1 i_0_85 (.A1(n_0_359), .A2(n_0_110), .B1(n_0_360), .B2(n_0_105), 
      .ZN(n_0_104));
   XOR2_X1 i_0_86 (.A(n_0_516), .B(n_0_106), .Z(n_0_105));
   NAND2_X1 i_0_87 (.A1(n_0_515), .A2(n_0_107), .ZN(n_0_106));
   AOI21_X1 i_0_88 (.A(in_e[1]), .B1(in_m[6]), .B2(n_0_109), .ZN(n_0_107));
   INV_X1 i_0_89 (.A(n_0_109), .ZN(n_0_108));
   AOI21_X1 i_0_90 (.A(n_0_157), .B1(in_e[1]), .B2(in_e[0]), .ZN(n_0_109));
   AOI221_X1 i_0_91 (.A(n_0_111), .B1(n_0_496), .B2(n_0_495), .C1(n_0_516), 
      .C2(n_0_112), .ZN(n_0_110));
   NOR2_X1 i_0_92 (.A1(n_0_516), .A2(n_0_112), .ZN(n_0_111));
   AOI21_X1 i_0_93 (.A(n_0_169), .B1(n_0_515), .B2(n_0_496), .ZN(n_0_112));
   INV_X1 i_0_94 (.A(n_0_114), .ZN(n_0_113));
   AOI21_X1 i_0_95 (.A(n_0_516), .B1(n_0_142), .B2(n_0_115), .ZN(n_0_114));
   AOI221_X1 i_0_96 (.A(n_0_177), .B1(n_0_464), .B2(n_0_22), .C1(n_0_12), 
      .C2(n_0_373), .ZN(n_0_115));
   NOR3_X1 i_0_97 (.A1(n_0_158), .A2(n_0_117), .A3(n_0_122), .ZN(n_0_116));
   AOI21_X1 i_0_98 (.A(n_0_121), .B1(n_0_484), .B2(n_0_118), .ZN(n_0_117));
   NAND3_X1 i_0_99 (.A1(n_0_495), .A2(n_0_198), .A3(n_0_119), .ZN(n_0_118));
   AOI221_X1 i_0_100 (.A(n_0_120), .B1(in_e[3]), .B2(in_m[15]), .C1(n_0_516), 
      .C2(in_m[7]), .ZN(n_0_119));
   NAND2_X1 i_0_101 (.A1(n_0_343), .A2(n_0_193), .ZN(n_0_120));
   AOI21_X1 i_0_102 (.A(n_0_156), .B1(in_e[3]), .B2(n_0_15), .ZN(n_0_121));
   NAND2_X1 i_0_103 (.A1(n_0_515), .A2(n_0_157), .ZN(n_0_15));
   NAND2_X1 i_0_104 (.A1(n_0_124), .A2(n_0_123), .ZN(n_0_122));
   AOI22_X1 i_0_105 (.A1(n_0_29), .A2(n_0_175), .B1(n_0_24), .B2(n_0_239), 
      .ZN(n_0_123));
   AOI221_X1 i_0_106 (.A(n_0_166), .B1(n_0_25), .B2(n_0_171), .C1(n_0_23), 
      .C2(n_0_261), .ZN(n_0_124));
   AOI222_X1 i_0_107 (.A1(n_0_26), .A2(n_0_164), .B1(n_0_28), .B2(n_0_179), 
      .C1(n_0_27), .C2(n_0_163), .ZN(n_0_125));
   INV_X1 i_0_108 (.A(n_0_126), .ZN(n_4));
   AOI221_X1 i_0_109 (.A(n_0_154), .B1(n_0_153), .B2(n_0_127), .C1(in_e[4]), 
      .C2(n_0_132), .ZN(n_0_126));
   NAND2_X1 i_0_110 (.A1(n_0_131), .A2(n_0_128), .ZN(n_0_127));
   AOI22_X1 i_0_111 (.A1(n_0_32), .A2(n_0_357), .B1(n_0_33), .B2(n_0_129), 
      .ZN(n_0_128));
   INV_X1 i_0_112 (.A(n_0_130), .ZN(n_0_129));
   NAND3_X1 i_0_113 (.A1(n_0_496), .A2(in_m[3]), .A3(n_0_359), .ZN(n_0_130));
   AOI22_X1 i_0_114 (.A1(n_0_31), .A2(n_0_151), .B1(in_m[6]), .B2(n_0_30), 
      .ZN(n_0_131));
   NAND4_X1 i_0_115 (.A1(n_0_139), .A2(n_0_137), .A3(n_0_133), .A4(n_0_140), 
      .ZN(n_0_132));
   AOI221_X1 i_0_116 (.A(n_0_134), .B1(n_0_0), .B2(n_0_171), .C1(n_0_188), 
      .C2(n_0_16), .ZN(n_0_133));
   INV_X1 i_0_117 (.A(n_0_135), .ZN(n_0_134));
   AOI221_X1 i_0_118 (.A(n_0_136), .B1(n_0_464), .B2(n_0_20), .C1(n_0_2), 
      .C2(n_0_261), .ZN(n_0_135));
   AOI21_X1 i_0_119 (.A(n_0_374), .B1(n_0_516), .B2(n_0_488), .ZN(n_0_136));
   AOI22_X1 i_0_120 (.A1(in_e[3]), .A2(n_0_138), .B1(n_0_1), .B2(n_0_239), 
      .ZN(n_0_137));
   NAND4_X1 i_0_121 (.A1(n_0_400), .A2(n_0_295), .A3(n_0_309), .A4(n_0_264), 
      .ZN(n_0_138));
   AOI22_X1 i_0_122 (.A1(n_0_4), .A2(n_0_163), .B1(n_0_6), .B2(n_0_175), 
      .ZN(n_0_139));
   AOI221_X1 i_0_123 (.A(n_0_141), .B1(n_0_5), .B2(n_0_179), .C1(n_0_3), 
      .C2(n_0_164), .ZN(n_0_140));
   INV_X1 i_0_124 (.A(n_0_142), .ZN(n_0_141));
   AOI221_X1 i_0_125 (.A(n_0_143), .B1(n_0_13), .B2(n_0_294), .C1(n_0_14), 
      .C2(n_0_308), .ZN(n_0_142));
   OAI22_X1 i_0_126 (.A1(n_0_514), .A2(n_0_404), .B1(n_0_515), .B2(n_0_400), 
      .ZN(n_0_143));
   INV_X1 i_0_127 (.A(n_0_144), .ZN(n_5));
   AOI21_X1 i_0_128 (.A(n_0_146), .B1(in_e[5]), .B2(n_0_147), .ZN(n_0_144));
   OAI21_X1 i_0_129 (.A(n_0_145), .B1(n_0_517), .B2(n_0_146), .ZN(n_6));
   XNOR2_X1 i_0_130 (.A(in_e[7]), .B(n_0_145), .ZN(n_7));
   NAND2_X1 i_0_131 (.A1(n_0_517), .A2(n_0_146), .ZN(n_0_145));
   NOR2_X1 i_0_132 (.A1(in_e[5]), .A2(n_0_147), .ZN(n_0_146));
   AOI21_X1 i_0_133 (.A(n_0_154), .B1(n_0_153), .B2(n_0_148), .ZN(n_0_147));
   OAI21_X1 i_0_134 (.A(n_0_149), .B1(n_0_9), .B2(n_0_358), .ZN(n_0_148));
   INV_X1 i_0_135 (.A(n_0_150), .ZN(n_0_149));
   AOI222_X1 i_0_136 (.A1(in_m[6]), .A2(n_0_7), .B1(n_0_8), .B2(n_0_151), 
      .C1(n_0_359), .C2(n_0_152), .ZN(n_0_150));
   NOR2_X1 i_0_137 (.A1(in_m[6]), .A2(n_0_497), .ZN(n_0_151));
   OR3_X1 i_0_138 (.A1(in_m[4]), .A2(n_0_495), .A3(n_0_10), .ZN(n_0_152));
   AND2_X1 i_0_139 (.A1(n_0_499), .A2(n_0_178), .ZN(n_0_153));
   AOI21_X1 i_0_140 (.A(in_e[4]), .B1(n_0_173), .B2(n_0_155), .ZN(n_0_154));
   AOI211_X1 i_0_141 (.A(n_0_158), .B(n_0_161), .C1(n_0_188), .C2(n_0_156), 
      .ZN(n_0_155));
   INV_X1 i_0_142 (.A(n_0_16), .ZN(n_0_156));
   NAND2_X1 i_0_143 (.A1(n_0_168), .A2(n_0_157), .ZN(n_0_16));
   INV_X1 i_0_144 (.A(n_0_157), .ZN(n_0_17));
   NOR2_X1 i_0_145 (.A1(in_e[1]), .A2(in_e[0]), .ZN(n_0_157));
   AOI21_X1 i_0_146 (.A(in_e[3]), .B1(n_0_160), .B2(n_0_159), .ZN(n_0_158));
   AOI221_X1 i_0_147 (.A(n_0_263), .B1(n_0_515), .B2(n_0_401), .C1(n_0_486), 
      .C2(n_0_294), .ZN(n_0_159));
   OR2_X1 i_0_148 (.A1(n_0_14), .A2(n_0_309), .ZN(n_0_160));
   OAI211_X1 i_0_149 (.A(n_0_165), .B(n_0_162), .C1(n_0_0), .C2(n_0_170), 
      .ZN(n_0_161));
   AOI22_X1 i_0_150 (.A1(n_0_490), .A2(n_0_164), .B1(n_0_489), .B2(n_0_163), 
      .ZN(n_0_162));
   AND2_X1 i_0_151 (.A1(in_m[10]), .A2(n_0_180), .ZN(n_0_163));
   NOR4_X1 i_0_152 (.A1(n_0_195), .A2(n_0_192), .A3(n_0_503), .A4(n_0_182), 
      .ZN(n_0_164));
   AOI21_X1 i_0_153 (.A(n_0_166), .B1(n_0_491), .B2(n_0_261), .ZN(n_0_165));
   OAI221_X1 i_0_154 (.A(n_0_167), .B1(n_0_404), .B2(n_0_18), .C1(n_0_465), 
      .C2(n_0_20), .ZN(n_0_166));
   NAND2_X1 i_0_155 (.A1(n_0_514), .A2(n_0_168), .ZN(n_0_18));
   NAND2_X1 i_0_156 (.A1(n_0_515), .A2(n_0_514), .ZN(n_0_19));
   NAND3_X1 i_0_157 (.A1(n_0_516), .A2(n_0_488), .A3(n_0_373), .ZN(n_0_167));
   NAND2_X1 i_0_158 (.A1(n_0_485), .A2(n_0_168), .ZN(n_0_20));
   INV_X1 i_0_159 (.A(n_0_21), .ZN(n_0_168));
   NAND2_X1 i_0_160 (.A1(n_0_516), .A2(n_0_515), .ZN(n_0_21));
   INV_X1 i_0_161 (.A(n_0_22), .ZN(n_0_169));
   NAND2_X1 i_0_162 (.A1(n_0_515), .A2(n_0_485), .ZN(n_0_22));
   INV_X1 i_0_163 (.A(n_0_171), .ZN(n_0_170));
   NOR3_X1 i_0_164 (.A1(n_0_195), .A2(n_0_192), .A3(n_0_172), .ZN(n_0_171));
   NAND2_X1 i_0_165 (.A1(in_m[12]), .A2(n_0_183), .ZN(n_0_172));
   AOI211_X1 i_0_166 (.A(n_0_177), .B(n_0_174), .C1(n_0_487), .C2(n_0_179), 
      .ZN(n_0_173));
   OAI22_X1 i_0_167 (.A1(n_0_6), .A2(n_0_176), .B1(n_0_1), .B2(n_0_238), 
      .ZN(n_0_174));
   INV_X1 i_0_168 (.A(n_0_176), .ZN(n_0_175));
   NAND2_X1 i_0_169 (.A1(n_0_281), .A2(n_0_180), .ZN(n_0_176));
   AND2_X1 i_0_170 (.A1(in_m[7]), .A2(n_0_178), .ZN(n_0_177));
   AND2_X1 i_0_171 (.A1(n_0_343), .A2(n_0_180), .ZN(n_0_178));
   AND2_X1 i_0_172 (.A1(n_0_311), .A2(n_0_180), .ZN(n_0_179));
   AND2_X1 i_0_173 (.A1(n_0_191), .A2(n_0_181), .ZN(n_0_180));
   INV_X1 i_0_174 (.A(n_0_182), .ZN(n_0_181));
   NAND2_X1 i_0_175 (.A1(n_0_504), .A2(n_0_183), .ZN(n_0_182));
   AND2_X1 i_0_176 (.A1(n_0_479), .A2(n_0_200), .ZN(n_0_183));
   AOI21_X1 i_0_177 (.A(in_m[23]), .B1(n_0_185), .B2(n_0_184), .ZN(n_8));
   NOR3_X1 i_0_178 (.A1(in_m[22]), .A2(n_0_433), .A3(n_0_254), .ZN(n_0_184));
   NOR3_X1 i_0_179 (.A1(in_m[9]), .A2(in_m[5]), .A3(n_0_186), .ZN(n_0_185));
   NAND3_X1 i_0_180 (.A1(n_0_512), .A2(n_0_428), .A3(n_0_187), .ZN(n_0_186));
   NOR4_X1 i_0_181 (.A1(in_m[10]), .A2(in_m[8]), .A3(in_m[4]), .A4(in_m[3]), 
      .ZN(n_0_187));
   NOR2_X1 i_0_182 (.A1(n_0_492), .A2(n_0_189), .ZN(n_9));
   OAI22_X1 i_0_183 (.A1(n_0_493), .A2(n_0_189), .B1(n_0_492), .B2(n_0_404), 
      .ZN(n_10));
   OAI222_X1 i_0_184 (.A1(n_0_492), .A2(n_0_465), .B1(n_0_493), .B2(n_0_404), 
      .C1(n_0_494), .C2(n_0_189), .ZN(n_11));
   INV_X1 i_0_185 (.A(n_0_189), .ZN(n_0_188));
   AOI21_X1 i_0_186 (.A(n_0_483), .B1(n_0_196), .B2(n_0_190), .ZN(n_0_189));
   AND3_X1 i_0_187 (.A1(n_0_499), .A2(n_0_495), .A3(n_0_191), .ZN(n_0_190));
   AND2_X1 i_0_188 (.A1(n_0_507), .A2(n_0_193), .ZN(n_0_191));
   NAND2_X1 i_0_189 (.A1(n_0_511), .A2(n_0_507), .ZN(n_0_192));
   NOR3_X1 i_0_190 (.A1(in_m[19]), .A2(in_m[11]), .A3(n_0_195), .ZN(n_0_193));
   INV_X1 i_0_191 (.A(n_0_195), .ZN(n_0_194));
   NAND2_X1 i_0_192 (.A1(n_0_505), .A2(n_0_476), .ZN(n_0_195));
   INV_X1 i_0_193 (.A(n_0_197), .ZN(n_0_196));
   NAND2_X1 i_0_194 (.A1(n_0_343), .A2(n_0_198), .ZN(n_0_197));
   NOR3_X1 i_0_195 (.A1(in_m[20]), .A2(in_m[4]), .A3(n_0_199), .ZN(n_0_198));
   NAND3_X1 i_0_196 (.A1(n_0_504), .A2(n_0_359), .A3(n_0_200), .ZN(n_0_199));
   NOR3_X1 i_0_197 (.A1(in_m[18]), .A2(in_m[16]), .A3(in_m[14]), .ZN(n_0_200));
   OAI221_X1 i_0_198 (.A(n_0_201), .B1(n_0_492), .B2(n_0_402), .C1(n_0_493), 
      .C2(n_0_465), .ZN(n_12));
   AOI22_X1 i_0_199 (.A1(in_m[2]), .A2(n_0_403), .B1(in_m[3]), .B2(n_0_483), 
      .ZN(n_0_201));
   OAI221_X1 i_0_200 (.A(n_0_202), .B1(n_0_493), .B2(n_0_402), .C1(n_0_494), 
      .C2(n_0_465), .ZN(n_13));
   AOI222_X1 i_0_201 (.A1(in_m[3]), .A2(n_0_403), .B1(in_m[4]), .B2(n_0_483), 
      .C1(in_m[0]), .C2(n_0_373), .ZN(n_0_202));
   OAI211_X1 i_0_202 (.A(n_0_204), .B(n_0_203), .C1(n_0_492), .C2(n_0_295), 
      .ZN(n_14));
   AOI22_X1 i_0_203 (.A1(in_m[1]), .A2(n_0_373), .B1(in_m[2]), .B2(n_0_401), 
      .ZN(n_0_203));
   AOI222_X1 i_0_204 (.A1(in_m[4]), .A2(n_0_403), .B1(in_m[5]), .B2(n_0_483), 
      .C1(in_m[3]), .C2(n_0_464), .ZN(n_0_204));
   OAI211_X1 i_0_205 (.A(n_0_205), .B(n_0_206), .C1(n_0_492), .C2(n_0_309), 
      .ZN(n_15));
   AOI222_X1 i_0_206 (.A1(in_m[5]), .A2(n_0_403), .B1(in_m[6]), .B2(n_0_483), 
      .C1(in_m[2]), .C2(n_0_373), .ZN(n_0_205));
   AOI222_X1 i_0_207 (.A1(in_m[1]), .A2(n_0_294), .B1(in_m[3]), .B2(n_0_401), 
      .C1(in_m[4]), .C2(n_0_464), .ZN(n_0_206));
   OAI211_X1 i_0_208 (.A(n_0_207), .B(n_0_209), .C1(n_0_493), .C2(n_0_309), 
      .ZN(n_16));
   AOI21_X1 i_0_209 (.A(n_0_208), .B1(in_m[0]), .B2(n_0_263), .ZN(n_0_207));
   OAI222_X1 i_0_210 (.A1(n_0_499), .A2(n_0_484), .B1(n_0_498), .B2(n_0_404), 
      .C1(n_0_497), .C2(n_0_465), .ZN(n_0_208));
   AOI222_X1 i_0_211 (.A1(in_m[3]), .A2(n_0_373), .B1(in_m[2]), .B2(n_0_294), 
      .C1(in_m[4]), .C2(n_0_401), .ZN(n_0_209));
   NAND4_X1 i_0_212 (.A1(n_0_214), .A2(n_0_212), .A3(n_0_211), .A4(n_0_210), 
      .ZN(n_17));
   NAND2_X1 i_0_213 (.A1(in_m[0]), .A2(n_0_261), .ZN(n_0_210));
   AOI222_X1 i_0_214 (.A1(in_m[6]), .A2(n_0_464), .B1(in_m[5]), .B2(n_0_401), 
      .C1(in_m[3]), .C2(n_0_294), .ZN(n_0_211));
   AOI221_X1 i_0_215 (.A(n_0_213), .B1(in_m[4]), .B2(n_0_373), .C1(in_m[1]), 
      .C2(n_0_263), .ZN(n_0_212));
   OAI22_X1 i_0_216 (.A1(n_0_499), .A2(n_0_404), .B1(n_0_500), .B2(n_0_484), 
      .ZN(n_0_213));
   NAND2_X1 i_0_217 (.A1(in_m[2]), .A2(n_0_308), .ZN(n_0_214));
   NAND4_X1 i_0_218 (.A1(n_0_219), .A2(n_0_217), .A3(n_0_215), .A4(n_0_220), 
      .ZN(n_18));
   AOI221_X1 i_0_219 (.A(n_0_216), .B1(in_m[5]), .B2(n_0_373), .C1(in_m[1]), 
      .C2(n_0_261), .ZN(n_0_215));
   OAI22_X1 i_0_220 (.A1(n_0_499), .A2(n_0_465), .B1(n_0_498), .B2(n_0_402), 
      .ZN(n_0_216));
   AOI21_X1 i_0_221 (.A(n_0_218), .B1(in_m[3]), .B2(n_0_308), .ZN(n_0_217));
   OAI222_X1 i_0_222 (.A1(n_0_500), .A2(n_0_404), .B1(n_0_501), .B2(n_0_484), 
      .C1(n_0_496), .C2(n_0_295), .ZN(n_0_218));
   NAND2_X1 i_0_223 (.A1(in_m[2]), .A2(n_0_263), .ZN(n_0_219));
   NAND2_X1 i_0_224 (.A1(in_m[0]), .A2(n_0_239), .ZN(n_0_220));
   NAND3_X1 i_0_225 (.A1(n_0_226), .A2(n_0_224), .A3(n_0_221), .ZN(n_19));
   AOI221_X1 i_0_226 (.A(n_0_222), .B1(in_m[3]), .B2(n_0_263), .C1(in_m[1]), 
      .C2(n_0_239), .ZN(n_0_221));
   OAI221_X1 i_0_227 (.A(n_0_223), .B1(n_0_499), .B2(n_0_402), .C1(n_0_496), 
      .C2(n_0_309), .ZN(n_0_222));
   AOI22_X1 i_0_228 (.A1(in_m[10]), .A2(n_0_483), .B1(in_m[9]), .B2(n_0_403), 
      .ZN(n_0_223));
   AOI221_X1 i_0_229 (.A(n_0_225), .B1(in_m[8]), .B2(n_0_464), .C1(in_m[2]), 
      .C2(n_0_261), .ZN(n_0_224));
   OAI22_X1 i_0_230 (.A1(n_0_498), .A2(n_0_374), .B1(n_0_497), .B2(n_0_295), 
      .ZN(n_0_225));
   NAND2_X1 i_0_231 (.A1(in_m[0]), .A2(n_0_233), .ZN(n_0_226));
   NAND4_X1 i_0_232 (.A1(n_0_228), .A2(n_0_227), .A3(n_0_231), .A4(n_0_232), 
      .ZN(n_20));
   AOI22_X1 i_0_233 (.A1(in_m[5]), .A2(n_0_308), .B1(in_m[4]), .B2(n_0_263), 
      .ZN(n_0_227));
   AOI211_X1 i_0_234 (.A(n_0_230), .B(n_0_229), .C1(in_m[6]), .C2(n_0_294), 
      .ZN(n_0_228));
   NOR3_X1 i_0_235 (.A1(n_0_492), .A2(n_0_319), .A3(n_0_254), .ZN(n_0_229));
   OAI22_X1 i_0_236 (.A1(n_0_503), .A2(n_0_484), .B1(n_0_502), .B2(n_0_404), 
      .ZN(n_0_230));
   NAND2_X1 i_0_237 (.A1(in_m[2]), .A2(n_0_239), .ZN(n_0_231));
   AOI221_X1 i_0_238 (.A(n_0_234), .B1(in_m[3]), .B2(n_0_261), .C1(in_m[1]), 
      .C2(n_0_233), .ZN(n_0_232));
   NOR2_X1 i_0_239 (.A1(n_0_451), .A2(n_0_368), .ZN(n_0_233));
   OAI222_X1 i_0_240 (.A1(n_0_500), .A2(n_0_402), .B1(n_0_499), .B2(n_0_374), 
      .C1(n_0_501), .C2(n_0_465), .ZN(n_0_234));
   OAI211_X1 i_0_241 (.A(n_0_235), .B(n_0_240), .C1(n_0_495), .C2(n_0_238), 
      .ZN(n_21));
   AOI211_X1 i_0_242 (.A(n_0_237), .B(n_0_236), .C1(in_m[6]), .C2(n_0_308), 
      .ZN(n_0_235));
   OAI33_X1 i_0_243 (.A1(n_0_492), .A2(n_0_310), .A3(n_0_292), .B1(n_0_494), 
      .B2(n_0_368), .B3(n_0_254), .ZN(n_0_236));
   NOR3_X1 i_0_244 (.A1(n_0_493), .A2(n_0_283), .A3(n_0_319), .ZN(n_0_237));
   INV_X1 i_0_245 (.A(n_0_239), .ZN(n_0_238));
   NOR3_X1 i_0_246 (.A1(n_0_394), .A2(n_0_254), .A3(n_0_483), .ZN(n_0_239));
   AOI211_X1 i_0_247 (.A(n_0_243), .B(n_0_241), .C1(in_m[4]), .C2(n_0_261), 
      .ZN(n_0_240));
   OAI221_X1 i_0_248 (.A(n_0_242), .B1(n_0_501), .B2(n_0_402), .C1(n_0_497), 
      .C2(n_0_264), .ZN(n_0_241));
   AOI22_X1 i_0_249 (.A1(in_m[12]), .A2(n_0_483), .B1(in_m[11]), .B2(n_0_403), 
      .ZN(n_0_242));
   OAI222_X1 i_0_250 (.A1(n_0_500), .A2(n_0_374), .B1(n_0_499), .B2(n_0_295), 
      .C1(n_0_502), .C2(n_0_465), .ZN(n_0_243));
   NAND4_X1 i_0_251 (.A1(n_0_246), .A2(n_0_244), .A3(n_0_248), .A4(n_0_251), 
      .ZN(n_22));
   INV_X1 i_0_252 (.A(n_0_245), .ZN(n_0_244));
   OAI33_X1 i_0_253 (.A1(n_0_495), .A2(n_0_368), .A3(n_0_283), .B1(n_0_494), 
      .B2(n_0_319), .B3(n_0_292), .ZN(n_0_245));
   AOI221_X1 i_0_254 (.A(n_0_247), .B1(in_m[9]), .B2(n_0_373), .C1(in_m[7]), 
      .C2(n_0_308), .ZN(n_0_246));
   OAI22_X1 i_0_255 (.A1(n_0_504), .A2(n_0_404), .B1(n_0_505), .B2(n_0_484), 
      .ZN(n_0_247));
   AOI211_X1 i_0_256 (.A(n_0_249), .B(n_0_250), .C1(in_m[6]), .C2(n_0_263), 
      .ZN(n_0_248));
   NOR3_X1 i_0_257 (.A1(n_0_493), .A2(n_0_310), .A3(n_0_314), .ZN(n_0_249));
   NOR3_X1 i_0_258 (.A1(n_0_492), .A2(n_0_297), .A3(n_0_348), .ZN(n_0_250));
   AOI211_X1 i_0_259 (.A(n_0_252), .B(n_0_253), .C1(in_m[5]), .C2(n_0_261), 
      .ZN(n_0_251));
   OAI222_X1 i_0_260 (.A1(n_0_503), .A2(n_0_465), .B1(n_0_500), .B2(n_0_295), 
      .C1(n_0_502), .C2(n_0_402), .ZN(n_0_252));
   NOR3_X1 i_0_261 (.A1(n_0_394), .A2(n_0_254), .A3(n_0_496), .ZN(n_0_253));
   NAND2_X1 i_0_262 (.A1(n_0_481), .A2(n_0_453), .ZN(n_0_254));
   NAND4_X1 i_0_263 (.A1(n_0_266), .A2(n_0_262), .A3(n_0_259), .A4(n_0_255), 
      .ZN(n_23));
   AOI211_X1 i_0_264 (.A(n_0_257), .B(n_0_256), .C1(in_m[13]), .C2(n_0_258), 
      .ZN(n_0_255));
   OAI33_X1 i_0_265 (.A1(n_0_494), .A2(n_0_310), .A3(n_0_348), .B1(n_0_495), 
      .B2(n_0_319), .B3(n_0_314), .ZN(n_0_256));
   OAI33_X1 i_0_266 (.A1(n_0_496), .A2(n_0_368), .A3(n_0_292), .B1(n_0_493), 
      .B2(n_0_297), .B3(n_0_364), .ZN(n_0_257));
   OAI33_X1 i_0_267 (.A1(in_m[23]), .A2(in_m[22]), .A3(n_0_513), .B1(in_m[14]), 
      .B2(n_0_497), .B3(n_0_283), .ZN(n_0_258));
   AOI221_X1 i_0_268 (.A(n_0_260), .B1(in_m[11]), .B2(n_0_401), .C1(in_m[6]), 
      .C2(n_0_261), .ZN(n_0_259));
   OAI22_X1 i_0_269 (.A1(n_0_501), .A2(n_0_295), .B1(n_0_502), .B2(n_0_374), 
      .ZN(n_0_260));
   NOR2_X1 i_0_270 (.A1(n_0_506), .A2(n_0_451), .ZN(n_0_261));
   AOI21_X1 i_0_271 (.A(n_0_265), .B1(in_m[7]), .B2(n_0_263), .ZN(n_0_262));
   INV_X1 i_0_272 (.A(n_0_264), .ZN(n_0_263));
   NAND2_X1 i_0_273 (.A1(n_0_477), .A2(n_0_322), .ZN(n_0_264));
   NOR3_X1 i_0_274 (.A1(n_0_492), .A2(n_0_280), .A3(n_0_367), .ZN(n_0_265));
   AOI222_X1 i_0_275 (.A1(in_m[12]), .A2(n_0_464), .B1(in_m[14]), .B2(n_0_483), 
      .C1(in_m[8]), .C2(n_0_308), .ZN(n_0_266));
   NAND4_X1 i_0_276 (.A1(n_0_268), .A2(n_0_267), .A3(n_0_275), .A4(n_0_270), 
      .ZN(n_24));
   AOI22_X1 i_0_277 (.A1(in_m[9]), .A2(n_0_308), .B1(in_m[14]), .B2(n_0_274), 
      .ZN(n_0_267));
   INV_X1 i_0_278 (.A(n_0_269), .ZN(n_0_268));
   OAI33_X1 i_0_279 (.A1(n_0_368), .A2(n_0_314), .A3(n_0_497), .B1(n_0_394), 
      .B2(n_0_292), .B3(n_0_498), .ZN(n_0_269));
   AND4_X1 i_0_280 (.A1(n_0_272), .A2(n_0_271), .A3(n_0_279), .A4(n_0_276), 
      .ZN(n_0_270));
   AOI221_X1 i_0_281 (.A(n_0_282), .B1(in_m[12]), .B2(n_0_401), .C1(in_m[15]), 
      .C2(n_0_483), .ZN(n_0_271));
   INV_X1 i_0_282 (.A(n_0_273), .ZN(n_0_272));
   OAI33_X1 i_0_283 (.A1(n_0_397), .A2(n_0_280), .A3(n_0_493), .B1(n_0_364), 
      .B2(n_0_310), .B3(n_0_495), .ZN(n_0_273));
   OAI21_X1 i_0_284 (.A(n_0_404), .B1(n_0_499), .B2(n_0_283), .ZN(n_0_274));
   NAND4_X1 i_0_285 (.A1(in_m[0]), .A2(n_0_338), .A3(in_m[7]), .A4(n_0_341), 
      .ZN(n_0_275));
   AOI221_X1 i_0_286 (.A(n_0_277), .B1(in_m[13]), .B2(n_0_464), .C1(in_m[11]), 
      .C2(n_0_373), .ZN(n_0_276));
   OAI21_X1 i_0_287 (.A(n_0_278), .B1(n_0_502), .B2(n_0_295), .ZN(n_0_277));
   NAND3_X1 i_0_288 (.A1(in_m[8]), .A2(n_0_481), .A3(n_0_322), .ZN(n_0_278));
   OR3_X1 i_0_289 (.A1(n_0_494), .A2(n_0_297), .A3(n_0_367), .ZN(n_0_279));
   NAND2_X1 i_0_290 (.A1(n_0_432), .A2(n_0_281), .ZN(n_0_280));
   NOR2_X1 i_0_291 (.A1(n_0_500), .A2(n_0_438), .ZN(n_0_281));
   NOR3_X1 i_0_292 (.A1(n_0_496), .A2(n_0_319), .A3(n_0_348), .ZN(n_0_282));
   NAND2_X1 i_0_293 (.A1(n_0_479), .A2(n_0_453), .ZN(n_0_283));
   NAND2_X1 i_0_294 (.A1(n_0_289), .A2(n_0_284), .ZN(n_25));
   NOR4_X1 i_0_295 (.A1(n_0_296), .A2(n_0_286), .A3(n_0_288), .A4(n_0_285), 
      .ZN(n_0_284));
   OAI33_X1 i_0_296 (.A1(n_0_364), .A2(n_0_319), .A3(n_0_497), .B1(n_0_394), 
      .B2(n_0_314), .B3(n_0_499), .ZN(n_0_285));
   OAI221_X1 i_0_297 (.A(n_0_287), .B1(n_0_507), .B2(n_0_404), .C1(n_0_504), 
      .C2(n_0_374), .ZN(n_0_286));
   AOI222_X1 i_0_298 (.A1(in_m[11]), .A2(n_0_294), .B1(n_0_455), .B2(n_0_290), 
      .C1(in_m[16]), .C2(n_0_483), .ZN(n_0_287));
   OAI33_X1 i_0_299 (.A1(n_0_511), .A2(n_0_478), .A3(n_0_505), .B1(n_0_368), 
      .B2(n_0_348), .B3(n_0_498), .ZN(n_0_288));
   AOI222_X1 i_0_300 (.A1(n_0_341), .A2(n_0_298), .B1(in_m[14]), .B2(n_0_291), 
      .C1(n_0_422), .C2(n_0_293), .ZN(n_0_289));
   OAI33_X1 i_0_301 (.A1(n_0_508), .A2(n_0_482), .A3(n_0_502), .B1(n_0_501), 
      .B2(n_0_372), .B3(n_0_480), .ZN(n_0_290));
   OAI21_X1 i_0_302 (.A(n_0_465), .B1(n_0_500), .B2(n_0_292), .ZN(n_0_291));
   NAND2_X1 i_0_303 (.A1(n_0_471), .A2(n_0_453), .ZN(n_0_292));
   NOR4_X1 i_0_304 (.A1(in_m[11]), .A2(n_0_494), .A3(n_0_500), .A4(n_0_421), 
      .ZN(n_0_293));
   INV_X1 i_0_305 (.A(n_0_295), .ZN(n_0_294));
   NAND2_X1 i_0_306 (.A1(n_0_477), .A2(n_0_365), .ZN(n_0_295));
   OAI33_X1 i_0_307 (.A1(n_0_495), .A2(n_0_297), .A3(n_0_397), .B1(n_0_496), 
      .B2(n_0_310), .B3(n_0_367), .ZN(n_0_296));
   NAND2_X1 i_0_308 (.A1(n_0_432), .A2(n_0_311), .ZN(n_0_297));
   OAI33_X1 i_0_309 (.A1(n_0_493), .A2(n_0_380), .A3(n_0_499), .B1(n_0_492), 
      .B2(n_0_445), .B3(n_0_417), .ZN(n_0_298));
   NAND4_X1 i_0_310 (.A1(n_0_305), .A2(n_0_303), .A3(n_0_301), .A4(n_0_299), 
      .ZN(n_26));
   AND4_X1 i_0_311 (.A1(n_0_321), .A2(n_0_320), .A3(n_0_307), .A4(n_0_300), 
      .ZN(n_0_299));
   NAND4_X1 i_0_312 (.A1(n_0_338), .A2(n_0_311), .A3(n_0_450), .A4(in_m[4]), 
      .ZN(n_0_300));
   AOI221_X1 i_0_313 (.A(n_0_302), .B1(in_m[14]), .B2(n_0_313), .C1(in_m[11]), 
      .C2(n_0_308), .ZN(n_0_301));
   NOR3_X1 i_0_314 (.A1(n_0_499), .A2(n_0_364), .A3(n_0_368), .ZN(n_0_302));
   AOI21_X1 i_0_315 (.A(n_0_304), .B1(in_m[8]), .B2(n_0_323), .ZN(n_0_303));
   OAI33_X1 i_0_316 (.A1(n_0_342), .A2(n_0_315), .A3(n_0_447), .B1(n_0_497), 
      .B2(n_0_346), .B3(n_0_356), .ZN(n_0_304));
   INV_X1 i_0_317 (.A(n_0_306), .ZN(n_0_305));
   OAI33_X1 i_0_318 (.A1(n_0_498), .A2(n_0_319), .A3(n_0_367), .B1(n_0_397), 
      .B2(n_0_310), .B3(n_0_497), .ZN(n_0_306));
   AOI21_X1 i_0_319 (.A(n_0_317), .B1(in_m[13]), .B2(n_0_373), .ZN(n_0_307));
   INV_X1 i_0_320 (.A(n_0_309), .ZN(n_0_308));
   NAND2_X1 i_0_321 (.A1(in_m[16]), .A2(n_0_454), .ZN(n_0_309));
   NAND2_X1 i_0_322 (.A1(in_m[10]), .A2(n_0_432), .ZN(n_0_310));
   INV_X1 i_0_323 (.A(n_0_312), .ZN(n_0_311));
   NAND2_X1 i_0_324 (.A1(n_0_502), .A2(in_m[9]), .ZN(n_0_312));
   OAI21_X1 i_0_325 (.A(n_0_402), .B1(n_0_501), .B2(n_0_314), .ZN(n_0_313));
   NAND3_X1 i_0_326 (.A1(n_0_510), .A2(n_0_509), .A3(n_0_452), .ZN(n_0_314));
   INV_X1 i_0_327 (.A(n_0_316), .ZN(n_0_315));
   OAI33_X1 i_0_328 (.A1(in_m[11]), .A2(n_0_494), .A3(n_0_499), .B1(in_m[12]), 
      .B2(n_0_417), .B3(n_0_493), .ZN(n_0_316));
   AOI21_X1 i_0_329 (.A(n_0_509), .B1(n_0_484), .B2(n_0_318), .ZN(n_0_317));
   NAND3_X1 i_0_330 (.A1(in_m[12]), .A2(n_0_467), .A3(n_0_481), .ZN(n_0_318));
   NAND2_X1 i_0_331 (.A1(in_m[11]), .A2(n_0_420), .ZN(n_0_319));
   NAND3_X1 i_0_332 (.A1(n_0_471), .A2(n_0_322), .A3(in_m[10]), .ZN(n_0_320));
   AOI22_X1 i_0_333 (.A1(in_m[16]), .A2(n_0_403), .B1(in_m[15]), .B2(n_0_464), 
      .ZN(n_0_321));
   NOR2_X1 i_0_334 (.A1(n_0_456), .A2(n_0_372), .ZN(n_0_322));
   OAI33_X1 i_0_335 (.A1(in_m[9]), .A2(n_0_495), .A3(n_0_333), .B1(in_m[14]), 
      .B2(n_0_505), .B3(n_0_348), .ZN(n_0_323));
   OAI211_X1 i_0_336 (.A(n_0_330), .B(n_0_324), .C1(n_0_356), .C2(n_0_349), 
      .ZN(n_27));
   NOR3_X1 i_0_337 (.A1(n_0_332), .A2(n_0_325), .A3(n_0_339), .ZN(n_0_324));
   INV_X1 i_0_338 (.A(n_0_326), .ZN(n_0_325));
   AOI211_X1 i_0_339 (.A(n_0_334), .B(n_0_327), .C1(in_m[18]), .C2(n_0_483), 
      .ZN(n_0_326));
   NAND3_X1 i_0_340 (.A1(n_0_337), .A2(n_0_328), .A3(n_0_329), .ZN(n_0_327));
   AOI221_X1 i_0_341 (.A(n_0_336), .B1(in_m[17]), .B2(n_0_403), .C1(n_0_470), 
      .C2(n_0_335), .ZN(n_0_328));
   NAND3_X1 i_0_342 (.A1(in_m[9]), .A2(n_0_363), .A3(n_0_393), .ZN(n_0_329));
   AOI21_X1 i_0_343 (.A(n_0_331), .B1(in_m[14]), .B2(n_0_347), .ZN(n_0_330));
   OAI33_X1 i_0_344 (.A1(n_0_368), .A2(n_0_367), .A3(n_0_500), .B1(n_0_496), 
      .B2(n_0_423), .B3(n_0_344), .ZN(n_0_331));
   AOI211_X1 i_0_345 (.A(n_0_497), .B(n_0_333), .C1(n_0_501), .C2(n_0_407), 
      .ZN(n_0_332));
   NAND3_X1 i_0_346 (.A1(n_0_502), .A2(n_0_379), .A3(n_0_450), .ZN(n_0_333));
   AOI21_X1 i_0_347 (.A(n_0_507), .B1(n_0_402), .B2(n_0_395), .ZN(n_0_334));
   OAI21_X1 i_0_348 (.A(n_0_512), .B1(n_0_504), .B2(n_0_456), .ZN(n_0_335));
   AND3_X1 i_0_349 (.A1(in_m[13]), .A2(n_0_479), .A3(n_0_365), .ZN(n_0_336));
   NAND4_X1 i_0_350 (.A1(in_m[10]), .A2(in_m[6]), .A3(n_0_338), .A4(n_0_450), 
      .ZN(n_0_337));
   NOR2_X1 i_0_351 (.A1(in_m[11]), .A2(n_0_421), .ZN(n_0_338));
   AOI211_X1 i_0_352 (.A(n_0_499), .B(n_0_419), .C1(n_0_395), .C2(n_0_340), 
      .ZN(n_0_339));
   NAND2_X1 i_0_353 (.A1(in_m[3]), .A2(n_0_341), .ZN(n_0_340));
   INV_X1 i_0_354 (.A(n_0_342), .ZN(n_0_341));
   NAND2_X1 i_0_355 (.A1(n_0_450), .A2(n_0_343), .ZN(n_0_342));
   NOR2_X1 i_0_356 (.A1(in_m[8]), .A2(n_0_438), .ZN(n_0_343));
   AOI21_X1 i_0_357 (.A(n_0_345), .B1(in_m[8]), .B2(n_0_444), .ZN(n_0_344));
   NOR3_X1 i_0_358 (.A1(in_m[5]), .A2(n_0_433), .A3(n_0_346), .ZN(n_0_345));
   NAND2_X1 i_0_359 (.A1(in_m[0]), .A2(n_0_428), .ZN(n_0_346));
   OAI22_X1 i_0_360 (.A1(n_0_482), .A2(n_0_376), .B1(n_0_502), .B2(n_0_348), 
      .ZN(n_0_347));
   NAND3_X1 i_0_361 (.A1(n_0_511), .A2(n_0_509), .A3(n_0_452), .ZN(n_0_348));
   NAND2_X1 i_0_362 (.A1(in_m[2]), .A2(n_0_416), .ZN(n_0_349));
   NAND4_X1 i_0_363 (.A1(n_0_354), .A2(n_0_352), .A3(n_0_377), .A4(n_0_350), 
      .ZN(n_28));
   INV_X1 i_0_364 (.A(n_0_351), .ZN(n_0_350));
   OAI33_X1 i_0_365 (.A1(n_0_496), .A2(n_0_356), .A3(n_0_499), .B1(n_0_394), 
      .B2(n_0_367), .B3(n_0_502), .ZN(n_0_351));
   AOI221_X1 i_0_366 (.A(n_0_353), .B1(in_m[19]), .B2(n_0_366), .C1(in_m[14]), 
      .C2(n_0_361), .ZN(n_0_352));
   NOR3_X1 i_0_367 (.A1(n_0_501), .A2(n_0_397), .A3(n_0_368), .ZN(n_0_353));
   AOI221_X1 i_0_368 (.A(n_0_369), .B1(in_m[17]), .B2(n_0_464), .C1(n_0_357), 
      .C2(n_0_355), .ZN(n_0_354));
   NOR3_X1 i_0_369 (.A1(n_0_493), .A2(n_0_431), .A3(n_0_423), .ZN(n_0_355));
   NAND3_X1 i_0_370 (.A1(n_0_501), .A2(n_0_450), .A3(n_0_430), .ZN(n_0_356));
   INV_X1 i_0_371 (.A(n_0_358), .ZN(n_0_357));
   NAND2_X1 i_0_372 (.A1(in_m[4]), .A2(n_0_359), .ZN(n_0_358));
   INV_X1 i_0_373 (.A(n_0_360), .ZN(n_0_359));
   NAND2_X1 i_0_374 (.A1(n_0_498), .A2(n_0_497), .ZN(n_0_360));
   INV_X1 i_0_375 (.A(n_0_362), .ZN(n_0_361));
   AOI22_X1 i_0_376 (.A1(n_0_471), .A2(n_0_365), .B1(in_m[11]), .B2(n_0_363), 
      .ZN(n_0_362));
   INV_X1 i_0_377 (.A(n_0_364), .ZN(n_0_363));
   NAND2_X1 i_0_378 (.A1(n_0_467), .A2(n_0_452), .ZN(n_0_364));
   NOR2_X1 i_0_379 (.A1(n_0_509), .A2(n_0_468), .ZN(n_0_365));
   OAI21_X1 i_0_380 (.A(n_0_484), .B1(n_0_508), .B2(n_0_478), .ZN(n_0_366));
   NAND2_X1 i_0_381 (.A1(n_0_507), .A2(n_0_454), .ZN(n_0_367));
   NAND2_X1 i_0_382 (.A1(in_m[12]), .A2(n_0_446), .ZN(n_0_368));
   OAI222_X1 i_0_383 (.A1(n_0_507), .A2(n_0_374), .B1(n_0_510), .B2(n_0_404), 
      .C1(n_0_475), .C2(n_0_370), .ZN(n_0_369));
   INV_X1 i_0_384 (.A(n_0_371), .ZN(n_0_370));
   OAI33_X1 i_0_385 (.A1(n_0_508), .A2(n_0_505), .A3(in_m[18]), .B1(in_m[19]), 
      .B2(n_0_372), .B3(n_0_504), .ZN(n_0_371));
   NAND2_X1 i_0_386 (.A1(n_0_508), .A2(in_m[15]), .ZN(n_0_372));
   INV_X1 i_0_387 (.A(n_0_374), .ZN(n_0_373));
   NAND2_X1 i_0_388 (.A1(n_0_477), .A2(n_0_375), .ZN(n_0_374));
   INV_X1 i_0_389 (.A(n_0_376), .ZN(n_0_375));
   NAND2_X1 i_0_390 (.A1(n_0_511), .A2(in_m[18]), .ZN(n_0_376));
   OAI21_X1 i_0_391 (.A(n_0_450), .B1(n_0_381), .B2(n_0_378), .ZN(n_0_377));
   OAI33_X1 i_0_392 (.A1(n_0_502), .A2(n_0_380), .A3(n_0_499), .B1(n_0_503), 
      .B2(n_0_421), .B3(n_0_500), .ZN(n_0_378));
   INV_X1 i_0_393 (.A(n_0_380), .ZN(n_0_379));
   NAND2_X1 i_0_394 (.A1(n_0_506), .A2(n_0_434), .ZN(n_0_380));
   AOI21_X1 i_0_395 (.A(in_m[10]), .B1(n_0_384), .B2(n_0_382), .ZN(n_0_381));
   OAI21_X1 i_0_396 (.A(n_0_383), .B1(in_m[6]), .B2(n_0_387), .ZN(n_0_382));
   OAI33_X1 i_0_397 (.A1(n_0_495), .A2(n_0_431), .A3(in_m[7]), .B1(n_0_501), 
      .B2(n_0_445), .B3(n_0_498), .ZN(n_0_383));
   NAND3_X1 i_0_398 (.A1(in_m[5]), .A2(n_0_385), .A3(n_0_501), .ZN(n_0_384));
   AOI21_X1 i_0_399 (.A(n_0_419), .B1(n_0_500), .B2(n_0_386), .ZN(n_0_385));
   NAND3_X1 i_0_400 (.A1(n_0_503), .A2(in_m[2]), .A3(n_0_428), .ZN(n_0_386));
   NOR4_X1 i_0_401 (.A1(in_m[9]), .A2(in_m[5]), .A3(in_m[4]), .A4(n_0_492), 
      .ZN(n_0_387));
   INV_X1 i_0_402 (.A(n_0_388), .ZN(n_29));
   AOI221_X1 i_0_403 (.A(n_0_390), .B1(n_0_507), .B2(n_0_389), .C1(n_0_450), 
      .C2(n_0_408), .ZN(n_0_388));
   OAI33_X1 i_0_404 (.A1(n_0_501), .A2(n_0_419), .A3(n_0_395), .B1(n_0_504), 
      .B2(n_0_456), .B3(n_0_473), .ZN(n_0_389));
   OAI221_X1 i_0_405 (.A(n_0_392), .B1(n_0_395), .B2(n_0_394), .C1(n_0_407), 
      .C2(n_0_391), .ZN(n_0_390));
   NAND3_X1 i_0_406 (.A1(n_0_496), .A2(in_m[3]), .A3(n_0_422), .ZN(n_0_391));
   NOR3_X1 i_0_407 (.A1(n_0_406), .A2(n_0_399), .A3(n_0_398), .ZN(n_0_392));
   INV_X1 i_0_408 (.A(n_0_394), .ZN(n_0_393));
   NAND2_X1 i_0_409 (.A1(n_0_506), .A2(in_m[13]), .ZN(n_0_394));
   NAND2_X1 i_0_410 (.A1(in_m[11]), .A2(n_0_396), .ZN(n_0_395));
   INV_X1 i_0_411 (.A(n_0_397), .ZN(n_0_396));
   NAND2_X1 i_0_412 (.A1(n_0_508), .A2(n_0_454), .ZN(n_0_397));
   AOI211_X1 i_0_413 (.A(in_m[19]), .B(n_0_508), .C1(n_0_473), .C2(n_0_466), 
      .ZN(n_0_398));
   OAI33_X1 i_0_414 (.A1(n_0_507), .A2(n_0_478), .A3(n_0_405), .B1(n_0_476), 
      .B2(n_0_400), .B3(n_0_511), .ZN(n_0_399));
   NOR2_X1 i_0_415 (.A1(n_0_403), .A2(n_0_401), .ZN(n_0_400));
   INV_X1 i_0_416 (.A(n_0_402), .ZN(n_0_401));
   NAND2_X1 i_0_417 (.A1(in_m[19]), .A2(n_0_477), .ZN(n_0_402));
   INV_X1 i_0_418 (.A(n_0_404), .ZN(n_0_403));
   NAND2_X1 i_0_419 (.A1(in_m[21]), .A2(n_0_484), .ZN(n_0_404));
   AOI21_X1 i_0_420 (.A(n_0_461), .B1(n_0_510), .B2(in_m[17]), .ZN(n_0_405));
   AOI21_X1 i_0_421 (.A(n_0_512), .B1(n_0_484), .B2(n_0_466), .ZN(n_0_406));
   NAND3_X1 i_0_422 (.A1(in_m[1]), .A2(n_0_430), .A3(n_0_428), .ZN(n_0_407));
   OAI21_X1 i_0_423 (.A(n_0_409), .B1(n_0_500), .B2(n_0_411), .ZN(n_0_408));
   AOI22_X1 i_0_424 (.A1(n_0_502), .A2(n_0_412), .B1(in_m[10]), .B2(n_0_410), 
      .ZN(n_0_409));
   OAI22_X1 i_0_425 (.A1(n_0_500), .A2(n_0_445), .B1(in_m[13]), .B2(n_0_504), 
      .ZN(n_0_410));
   NAND3_X1 i_0_426 (.A1(in_m[6]), .A2(n_0_432), .A3(n_0_501), .ZN(n_0_411));
   OAI33_X1 i_0_427 (.A1(n_0_416), .A2(n_0_415), .A3(n_0_418), .B1(in_m[9]), 
      .B2(n_0_413), .B3(n_0_436), .ZN(n_0_412));
   INV_X1 i_0_428 (.A(n_0_414), .ZN(n_0_413));
   OAI33_X1 i_0_429 (.A1(in_m[12]), .A2(n_0_445), .A3(n_0_498), .B1(in_m[5]), 
      .B2(n_0_494), .B3(n_0_431), .ZN(n_0_414));
   AOI21_X1 i_0_430 (.A(in_m[7]), .B1(n_0_501), .B2(in_m[3]), .ZN(n_0_415));
   INV_X1 i_0_431 (.A(n_0_417), .ZN(n_0_416));
   NAND2_X1 i_0_432 (.A1(n_0_499), .A2(in_m[6]), .ZN(n_0_417));
   AOI22_X1 i_0_433 (.A1(in_m[5]), .A2(n_0_430), .B1(in_m[9]), .B2(n_0_420), 
      .ZN(n_0_418));
   INV_X1 i_0_434 (.A(n_0_420), .ZN(n_0_419));
   NOR2_X1 i_0_435 (.A1(in_m[14]), .A2(n_0_421), .ZN(n_0_420));
   NAND2_X1 i_0_436 (.A1(n_0_505), .A2(n_0_504), .ZN(n_0_421));
   OAI211_X1 i_0_437 (.A(n_0_462), .B(n_0_457), .C1(n_0_451), .C2(n_0_424), 
      .ZN(n_30));
   INV_X1 i_0_438 (.A(n_0_423), .ZN(n_0_422));
   NAND2_X1 i_0_439 (.A1(n_0_450), .A2(n_0_437), .ZN(n_0_423));
   AOI21_X1 i_0_440 (.A(n_0_439), .B1(n_0_437), .B2(n_0_425), .ZN(n_0_424));
   OAI33_X1 i_0_441 (.A1(n_0_498), .A2(n_0_433), .A3(n_0_499), .B1(in_m[8]), 
      .B2(n_0_433), .B3(n_0_426), .ZN(n_0_425));
   AOI21_X1 i_0_442 (.A(n_0_427), .B1(in_m[5]), .B2(n_0_435), .ZN(n_0_426));
   AND3_X1 i_0_443 (.A1(in_m[3]), .A2(n_0_428), .A3(n_0_429), .ZN(n_0_427));
   NOR2_X1 i_0_444 (.A1(in_m[7]), .A2(in_m[6]), .ZN(n_0_428));
   OAI21_X1 i_0_445 (.A(n_0_496), .B1(in_m[5]), .B2(n_0_494), .ZN(n_0_429));
   INV_X1 i_0_446 (.A(n_0_431), .ZN(n_0_430));
   NAND2_X1 i_0_447 (.A1(n_0_500), .A2(n_0_432), .ZN(n_0_431));
   INV_X1 i_0_448 (.A(n_0_433), .ZN(n_0_432));
   NAND2_X1 i_0_449 (.A1(n_0_446), .A2(n_0_434), .ZN(n_0_433));
   NOR2_X1 i_0_450 (.A1(in_m[12]), .A2(in_m[11]), .ZN(n_0_434));
   NAND2_X1 i_0_451 (.A1(n_0_498), .A2(n_0_436), .ZN(n_0_435));
   NAND2_X1 i_0_452 (.A1(n_0_499), .A2(in_m[4]), .ZN(n_0_436));
   INV_X1 i_0_453 (.A(n_0_438), .ZN(n_0_437));
   NAND2_X1 i_0_454 (.A1(n_0_502), .A2(n_0_501), .ZN(n_0_438));
   AOI21_X1 i_0_455 (.A(n_0_443), .B1(n_0_503), .B2(n_0_440), .ZN(n_0_439));
   INV_X1 i_0_456 (.A(n_0_441), .ZN(n_0_440));
   AOI21_X1 i_0_457 (.A(n_0_442), .B1(n_0_505), .B2(in_m[12]), .ZN(n_0_441));
   AOI211_X1 i_0_458 (.A(in_m[12]), .B(in_m[9]), .C1(n_0_502), .C2(in_m[7]), 
      .ZN(n_0_442));
   AOI22_X1 i_0_459 (.A1(n_0_449), .A2(n_0_448), .B1(in_m[8]), .B2(n_0_444), 
      .ZN(n_0_443));
   INV_X1 i_0_460 (.A(n_0_445), .ZN(n_0_444));
   NAND2_X1 i_0_461 (.A1(n_0_503), .A2(n_0_446), .ZN(n_0_445));
   INV_X1 i_0_462 (.A(n_0_447), .ZN(n_0_446));
   NAND2_X1 i_0_463 (.A1(n_0_506), .A2(n_0_505), .ZN(n_0_447));
   NAND2_X1 i_0_464 (.A1(in_m[14]), .A2(n_0_505), .ZN(n_0_448));
   OAI21_X1 i_0_465 (.A(n_0_504), .B1(in_m[13]), .B2(n_0_502), .ZN(n_0_449));
   INV_X1 i_0_466 (.A(n_0_451), .ZN(n_0_450));
   NAND2_X1 i_0_467 (.A1(n_0_455), .A2(n_0_452), .ZN(n_0_451));
   NOR3_X1 i_0_468 (.A1(in_m[16]), .A2(in_m[15]), .A3(n_0_478), .ZN(n_0_452));
   NOR3_X1 i_0_469 (.A1(in_m[16]), .A2(in_m[15]), .A3(n_0_456), .ZN(n_0_453));
   NOR2_X1 i_0_470 (.A1(n_0_478), .A2(n_0_456), .ZN(n_0_454));
   INV_X1 i_0_471 (.A(n_0_456), .ZN(n_0_455));
   NAND2_X1 i_0_472 (.A1(n_0_509), .A2(n_0_467), .ZN(n_0_456));
   INV_X1 i_0_473 (.A(n_0_458), .ZN(n_0_457));
   OAI33_X1 i_0_474 (.A1(n_0_469), .A2(n_0_468), .A3(n_0_507), .B1(n_0_460), 
      .B2(n_0_459), .B3(n_0_478), .ZN(n_0_458));
   AOI211_X1 i_0_475 (.A(in_m[18]), .B(n_0_509), .C1(n_0_511), .C2(in_m[16]), 
      .ZN(n_0_459));
   AOI21_X1 i_0_476 (.A(in_m[17]), .B1(in_m[14]), .B2(n_0_461), .ZN(n_0_460));
   NOR3_X1 i_0_477 (.A1(in_m[16]), .A2(n_0_505), .A3(n_0_468), .ZN(n_0_461));
   AOI21_X1 i_0_478 (.A(n_0_463), .B1(in_m[21]), .B2(n_0_480), .ZN(n_0_462));
   AOI21_X1 i_0_479 (.A(n_0_511), .B1(n_0_466), .B2(n_0_465), .ZN(n_0_463));
   INV_X1 i_0_480 (.A(n_0_465), .ZN(n_0_464));
   NAND2_X1 i_0_481 (.A1(in_m[20]), .A2(n_0_471), .ZN(n_0_465));
   NAND2_X1 i_0_482 (.A1(in_m[18]), .A2(n_0_471), .ZN(n_0_466));
   INV_X1 i_0_483 (.A(n_0_468), .ZN(n_0_467));
   NAND2_X1 i_0_484 (.A1(n_0_511), .A2(n_0_510), .ZN(n_0_468));
   AOI21_X1 i_0_485 (.A(n_0_474), .B1(n_0_512), .B2(n_0_470), .ZN(n_0_469));
   NOR2_X1 i_0_486 (.A1(n_0_508), .A2(n_0_472), .ZN(n_0_470));
   INV_X1 i_0_487 (.A(n_0_472), .ZN(n_0_471));
   NAND2_X1 i_0_488 (.A1(n_0_513), .A2(n_0_484), .ZN(n_0_472));
   INV_X1 i_0_489 (.A(n_0_474), .ZN(n_0_473));
   NOR2_X1 i_0_490 (.A1(n_0_506), .A2(n_0_475), .ZN(n_0_474));
   NAND2_X1 i_0_491 (.A1(n_0_479), .A2(n_0_476), .ZN(n_0_475));
   NOR2_X1 i_0_492 (.A1(in_m[21]), .A2(in_m[17]), .ZN(n_0_476));
   INV_X1 i_0_493 (.A(n_0_478), .ZN(n_0_477));
   NAND2_X1 i_0_494 (.A1(n_0_513), .A2(n_0_479), .ZN(n_0_478));
   INV_X1 i_0_495 (.A(n_0_480), .ZN(n_0_479));
   NAND2_X1 i_0_496 (.A1(n_0_512), .A2(n_0_484), .ZN(n_0_480));
   INV_X1 i_0_497 (.A(n_0_482), .ZN(n_0_481));
   NAND2_X1 i_0_498 (.A1(n_0_513), .A2(n_0_512), .ZN(n_0_482));
   INV_X1 i_0_499 (.A(n_0_484), .ZN(n_0_483));
   NOR2_X1 i_0_500 (.A1(in_m[23]), .A2(in_m[22]), .ZN(n_0_484));
   INV_X1 i_0_501 (.A(n_0_11), .ZN(n_0_485));
   INV_X1 i_0_502 (.A(n_0_13), .ZN(n_0_486));
   INV_X1 i_0_503 (.A(n_0_5), .ZN(n_0_487));
   INV_X1 i_0_504 (.A(n_0_12), .ZN(n_0_488));
   INV_X1 i_0_505 (.A(n_0_4), .ZN(n_0_489));
   INV_X1 i_0_506 (.A(n_0_3), .ZN(n_0_490));
   INV_X1 i_0_507 (.A(n_0_2), .ZN(n_0_491));
   INV_X1 i_0_508 (.A(in_m[0]), .ZN(n_0_492));
   INV_X1 i_0_509 (.A(in_m[1]), .ZN(n_0_493));
   INV_X1 i_0_510 (.A(in_m[2]), .ZN(n_0_494));
   INV_X1 i_0_511 (.A(in_m[3]), .ZN(n_0_495));
   INV_X1 i_0_512 (.A(in_m[4]), .ZN(n_0_496));
   INV_X1 i_0_513 (.A(in_m[5]), .ZN(n_0_497));
   INV_X1 i_0_514 (.A(in_m[6]), .ZN(n_0_498));
   INV_X1 i_0_515 (.A(in_m[7]), .ZN(n_0_499));
   INV_X1 i_0_516 (.A(in_m[8]), .ZN(n_0_500));
   INV_X1 i_0_517 (.A(in_m[9]), .ZN(n_0_501));
   INV_X1 i_0_518 (.A(in_m[10]), .ZN(n_0_502));
   INV_X1 i_0_519 (.A(in_m[11]), .ZN(n_0_503));
   INV_X1 i_0_520 (.A(in_m[12]), .ZN(n_0_504));
   INV_X1 i_0_521 (.A(in_m[13]), .ZN(n_0_505));
   INV_X1 i_0_522 (.A(in_m[14]), .ZN(n_0_506));
   INV_X1 i_0_523 (.A(in_m[15]), .ZN(n_0_507));
   INV_X1 i_0_524 (.A(in_m[16]), .ZN(n_0_508));
   INV_X1 i_0_525 (.A(in_m[17]), .ZN(n_0_509));
   INV_X1 i_0_526 (.A(in_m[18]), .ZN(n_0_510));
   INV_X1 i_0_527 (.A(in_m[19]), .ZN(n_0_511));
   INV_X1 i_0_528 (.A(in_m[20]), .ZN(n_0_512));
   INV_X1 i_0_529 (.A(in_m[21]), .ZN(n_0_513));
   INV_X1 i_0_530 (.A(in_e[1]), .ZN(n_0_514));
   INV_X1 i_0_531 (.A(in_e[2]), .ZN(n_0_515));
   INV_X1 i_0_532 (.A(in_e[3]), .ZN(n_0_516));
   INV_X1 i_0_533 (.A(in_e[6]), .ZN(n_0_517));
endmodule

module datapath__0_57(p_0, p_1, p_2);
   input [23:0]p_0;
   output [24:0]p_1;
   input [23:0]p_2;

   INV_X1 i_0 (.A(p_0[0]), .ZN(n_0));
   NAND2_X1 i_1 (.A1(n_0), .A2(p_2[0]), .ZN(n_1));
   OAI21_X1 i_2 (.A(n_1), .B1(p_2[0]), .B2(n_0), .ZN(p_1[0]));
   XNOR2_X1 i_3 (.A(p_0[1]), .B(p_2[1]), .ZN(n_2));
   XOR2_X1 i_4 (.A(n_2), .B(n_1), .Z(p_1[1]));
   INV_X1 i_5 (.A(n_1), .ZN(n_3));
   INV_X1 i_6 (.A(p_0[1]), .ZN(n_4));
   AOI22_X1 i_7 (.A1(n_2), .A2(n_3), .B1(n_4), .B2(p_2[1]), .ZN(n_5));
   XOR2_X1 i_8 (.A(p_0[2]), .B(p_2[2]), .Z(n_6));
   XNOR2_X1 i_9 (.A(n_5), .B(n_6), .ZN(p_1[2]));
   INV_X1 i_10 (.A(p_2[2]), .ZN(n_7));
   OAI22_X1 i_11 (.A1(n_5), .A2(n_6), .B1(n_7), .B2(p_0[2]), .ZN(n_8));
   XNOR2_X1 i_12 (.A(p_0[3]), .B(p_2[3]), .ZN(n_9));
   XNOR2_X1 i_13 (.A(n_8), .B(n_9), .ZN(p_1[3]));
   INV_X1 i_14 (.A(p_0[3]), .ZN(n_10));
   AOI22_X1 i_15 (.A1(n_8), .A2(n_9), .B1(n_10), .B2(p_2[3]), .ZN(n_11));
   XOR2_X1 i_16 (.A(p_0[4]), .B(p_2[4]), .Z(n_12));
   XNOR2_X1 i_17 (.A(n_11), .B(n_12), .ZN(p_1[4]));
   INV_X1 i_18 (.A(p_2[4]), .ZN(n_13));
   OAI22_X1 i_19 (.A1(n_11), .A2(n_12), .B1(n_13), .B2(p_0[4]), .ZN(n_14));
   XNOR2_X1 i_20 (.A(p_0[5]), .B(p_2[5]), .ZN(n_15));
   XNOR2_X1 i_21 (.A(n_14), .B(n_15), .ZN(p_1[5]));
   INV_X1 i_22 (.A(p_0[5]), .ZN(n_16));
   AOI22_X1 i_23 (.A1(n_14), .A2(n_15), .B1(n_16), .B2(p_2[5]), .ZN(n_17));
   XOR2_X1 i_24 (.A(p_0[6]), .B(p_2[6]), .Z(n_18));
   XNOR2_X1 i_25 (.A(n_17), .B(n_18), .ZN(p_1[6]));
   INV_X1 i_26 (.A(p_2[6]), .ZN(n_19));
   OAI22_X1 i_27 (.A1(n_17), .A2(n_18), .B1(n_19), .B2(p_0[6]), .ZN(n_20));
   XNOR2_X1 i_28 (.A(p_0[7]), .B(p_2[7]), .ZN(n_21));
   XNOR2_X1 i_29 (.A(n_20), .B(n_21), .ZN(p_1[7]));
   INV_X1 i_30 (.A(p_0[7]), .ZN(n_22));
   AOI22_X1 i_31 (.A1(n_20), .A2(n_21), .B1(n_22), .B2(p_2[7]), .ZN(n_23));
   XOR2_X1 i_32 (.A(p_0[8]), .B(p_2[8]), .Z(n_24));
   XNOR2_X1 i_33 (.A(n_23), .B(n_24), .ZN(p_1[8]));
   INV_X1 i_34 (.A(p_2[8]), .ZN(n_25));
   OAI22_X1 i_35 (.A1(n_23), .A2(n_24), .B1(n_25), .B2(p_0[8]), .ZN(n_26));
   XNOR2_X1 i_36 (.A(p_0[9]), .B(p_2[9]), .ZN(n_27));
   XNOR2_X1 i_37 (.A(n_26), .B(n_27), .ZN(p_1[9]));
   INV_X1 i_38 (.A(p_0[9]), .ZN(n_28));
   AOI22_X1 i_39 (.A1(n_26), .A2(n_27), .B1(n_28), .B2(p_2[9]), .ZN(n_29));
   XOR2_X1 i_40 (.A(p_0[10]), .B(p_2[10]), .Z(n_30));
   XNOR2_X1 i_41 (.A(n_29), .B(n_30), .ZN(p_1[10]));
   INV_X1 i_42 (.A(p_2[10]), .ZN(n_31));
   OAI22_X1 i_43 (.A1(n_29), .A2(n_30), .B1(n_31), .B2(p_0[10]), .ZN(n_32));
   XNOR2_X1 i_44 (.A(p_0[11]), .B(p_2[11]), .ZN(n_33));
   XNOR2_X1 i_45 (.A(n_32), .B(n_33), .ZN(p_1[11]));
   INV_X1 i_46 (.A(p_0[11]), .ZN(n_34));
   AOI22_X1 i_47 (.A1(n_32), .A2(n_33), .B1(n_34), .B2(p_2[11]), .ZN(n_35));
   XOR2_X1 i_48 (.A(p_0[12]), .B(p_2[12]), .Z(n_36));
   XNOR2_X1 i_49 (.A(n_35), .B(n_36), .ZN(p_1[12]));
   INV_X1 i_50 (.A(p_2[12]), .ZN(n_37));
   OAI22_X1 i_51 (.A1(n_35), .A2(n_36), .B1(n_37), .B2(p_0[12]), .ZN(n_38));
   XNOR2_X1 i_52 (.A(p_0[13]), .B(p_2[13]), .ZN(n_39));
   XNOR2_X1 i_53 (.A(n_38), .B(n_39), .ZN(p_1[13]));
   INV_X1 i_54 (.A(p_0[13]), .ZN(n_40));
   AOI22_X1 i_55 (.A1(n_38), .A2(n_39), .B1(n_40), .B2(p_2[13]), .ZN(n_41));
   INV_X1 i_56 (.A(n_41), .ZN(n_42));
   INV_X1 i_57 (.A(p_2[14]), .ZN(n_43));
   NAND2_X1 i_58 (.A1(n_43), .A2(p_0[14]), .ZN(n_44));
   INV_X1 i_59 (.A(n_44), .ZN(n_45));
   OR2_X1 i_60 (.A1(n_43), .A2(p_0[14]), .ZN(n_46));
   AOI21_X1 i_61 (.A(n_45), .B1(n_41), .B2(n_46), .ZN(n_47));
   NAND2_X1 i_62 (.A1(n_47), .A2(n_46), .ZN(n_48));
   INV_X1 i_63 (.A(n_47), .ZN(n_49));
   AOI22_X1 i_64 (.A1(n_42), .A2(n_48), .B1(n_49), .B2(n_44), .ZN(p_1[14]));
   XNOR2_X1 i_65 (.A(p_0[15]), .B(p_2[15]), .ZN(n_50));
   XNOR2_X1 i_66 (.A(n_47), .B(n_50), .ZN(p_1[15]));
   INV_X1 i_67 (.A(p_0[15]), .ZN(n_51));
   AOI22_X1 i_68 (.A1(n_47), .A2(n_50), .B1(n_51), .B2(p_2[15]), .ZN(n_52));
   XOR2_X1 i_69 (.A(p_0[16]), .B(p_2[16]), .Z(n_53));
   XNOR2_X1 i_70 (.A(n_52), .B(n_53), .ZN(p_1[16]));
   INV_X1 i_71 (.A(p_2[16]), .ZN(n_54));
   OAI22_X1 i_72 (.A1(n_52), .A2(n_53), .B1(n_54), .B2(p_0[16]), .ZN(n_55));
   XNOR2_X1 i_73 (.A(p_0[17]), .B(p_2[17]), .ZN(n_56));
   XNOR2_X1 i_74 (.A(n_55), .B(n_56), .ZN(p_1[17]));
   INV_X1 i_75 (.A(p_0[17]), .ZN(n_57));
   AOI22_X1 i_76 (.A1(n_55), .A2(n_56), .B1(n_57), .B2(p_2[17]), .ZN(n_58));
   XOR2_X1 i_77 (.A(p_0[18]), .B(p_2[18]), .Z(n_59));
   XNOR2_X1 i_78 (.A(n_58), .B(n_59), .ZN(p_1[18]));
   INV_X1 i_79 (.A(p_2[18]), .ZN(n_60));
   OAI22_X1 i_80 (.A1(n_58), .A2(n_59), .B1(n_60), .B2(p_0[18]), .ZN(n_61));
   XNOR2_X1 i_81 (.A(p_0[19]), .B(p_2[19]), .ZN(n_62));
   XNOR2_X1 i_82 (.A(n_61), .B(n_62), .ZN(p_1[19]));
   INV_X1 i_83 (.A(p_0[19]), .ZN(n_63));
   AOI22_X1 i_84 (.A1(n_61), .A2(n_62), .B1(n_63), .B2(p_2[19]), .ZN(n_64));
   INV_X1 i_85 (.A(n_64), .ZN(n_65));
   INV_X1 i_86 (.A(p_2[20]), .ZN(n_66));
   NAND2_X1 i_87 (.A1(n_66), .A2(p_0[20]), .ZN(n_67));
   INV_X1 i_88 (.A(n_67), .ZN(n_68));
   OR2_X1 i_89 (.A1(n_66), .A2(p_0[20]), .ZN(n_69));
   AOI21_X1 i_90 (.A(n_68), .B1(n_64), .B2(n_69), .ZN(n_70));
   NAND2_X1 i_91 (.A1(n_70), .A2(n_69), .ZN(n_71));
   INV_X1 i_92 (.A(n_70), .ZN(n_72));
   AOI22_X1 i_93 (.A1(n_65), .A2(n_71), .B1(n_72), .B2(n_67), .ZN(p_1[20]));
   XNOR2_X1 i_94 (.A(p_0[21]), .B(p_2[21]), .ZN(n_73));
   XNOR2_X1 i_95 (.A(n_70), .B(n_73), .ZN(p_1[21]));
   INV_X1 i_96 (.A(p_0[21]), .ZN(n_74));
   AOI22_X1 i_97 (.A1(n_70), .A2(n_73), .B1(n_74), .B2(p_2[21]), .ZN(n_75));
   XOR2_X1 i_98 (.A(p_0[22]), .B(p_2[22]), .Z(n_76));
   XNOR2_X1 i_99 (.A(n_75), .B(n_76), .ZN(p_1[22]));
   INV_X1 i_100 (.A(p_2[22]), .ZN(n_77));
   OAI22_X1 i_101 (.A1(n_75), .A2(n_76), .B1(n_77), .B2(p_0[22]), .ZN(n_78));
   XOR2_X1 i_102 (.A(p_2[23]), .B(p_0[23]), .Z(n_79));
   XOR2_X1 i_103 (.A(n_78), .B(n_79), .Z(p_1[23]));
   INV_X1 i_104 (.A(n_78), .ZN(n_80));
   INV_X1 i_105 (.A(p_2[23]), .ZN(n_81));
   OAI22_X1 i_106 (.A1(n_80), .A2(n_79), .B1(n_81), .B2(p_0[23]), .ZN(p_1[24]));
endmodule

module datapath__0_62(p_0, p_1, p_2);
   input [23:0]p_0;
   output [24:0]p_1;
   input [23:0]p_2;

   INV_X1 i_0 (.A(p_0[0]), .ZN(n_0));
   NAND2_X1 i_1 (.A1(n_0), .A2(p_2[0]), .ZN(n_1));
   OAI21_X1 i_2 (.A(n_1), .B1(p_2[0]), .B2(n_0), .ZN(p_1[0]));
   XNOR2_X1 i_3 (.A(p_0[1]), .B(p_2[1]), .ZN(n_2));
   XOR2_X1 i_4 (.A(n_2), .B(n_1), .Z(p_1[1]));
   INV_X1 i_5 (.A(n_1), .ZN(n_3));
   INV_X1 i_6 (.A(p_0[1]), .ZN(n_4));
   AOI22_X1 i_7 (.A1(n_2), .A2(n_3), .B1(n_4), .B2(p_2[1]), .ZN(n_5));
   XOR2_X1 i_8 (.A(p_0[2]), .B(p_2[2]), .Z(n_6));
   XNOR2_X1 i_9 (.A(n_5), .B(n_6), .ZN(p_1[2]));
   INV_X1 i_10 (.A(p_2[2]), .ZN(n_7));
   OAI22_X1 i_11 (.A1(n_5), .A2(n_6), .B1(n_7), .B2(p_0[2]), .ZN(n_8));
   XNOR2_X1 i_12 (.A(p_0[3]), .B(p_2[3]), .ZN(n_9));
   XNOR2_X1 i_13 (.A(n_8), .B(n_9), .ZN(p_1[3]));
   INV_X1 i_14 (.A(p_0[3]), .ZN(n_10));
   AOI22_X1 i_15 (.A1(n_8), .A2(n_9), .B1(n_10), .B2(p_2[3]), .ZN(n_11));
   XOR2_X1 i_16 (.A(p_0[4]), .B(p_2[4]), .Z(n_12));
   XNOR2_X1 i_17 (.A(n_11), .B(n_12), .ZN(p_1[4]));
   INV_X1 i_18 (.A(p_2[4]), .ZN(n_13));
   OAI22_X1 i_19 (.A1(n_11), .A2(n_12), .B1(n_13), .B2(p_0[4]), .ZN(n_14));
   XNOR2_X1 i_20 (.A(p_0[5]), .B(p_2[5]), .ZN(n_15));
   XNOR2_X1 i_21 (.A(n_14), .B(n_15), .ZN(p_1[5]));
   INV_X1 i_22 (.A(p_0[5]), .ZN(n_16));
   AOI22_X1 i_23 (.A1(n_14), .A2(n_15), .B1(n_16), .B2(p_2[5]), .ZN(n_17));
   XOR2_X1 i_24 (.A(p_0[6]), .B(p_2[6]), .Z(n_18));
   XNOR2_X1 i_25 (.A(n_17), .B(n_18), .ZN(p_1[6]));
   INV_X1 i_26 (.A(p_2[6]), .ZN(n_19));
   OAI22_X1 i_27 (.A1(n_17), .A2(n_18), .B1(n_19), .B2(p_0[6]), .ZN(n_20));
   XNOR2_X1 i_28 (.A(p_0[7]), .B(p_2[7]), .ZN(n_21));
   XNOR2_X1 i_29 (.A(n_20), .B(n_21), .ZN(p_1[7]));
   INV_X1 i_30 (.A(p_0[7]), .ZN(n_22));
   AOI22_X1 i_31 (.A1(n_20), .A2(n_21), .B1(n_22), .B2(p_2[7]), .ZN(n_23));
   XOR2_X1 i_32 (.A(p_0[8]), .B(p_2[8]), .Z(n_24));
   XNOR2_X1 i_33 (.A(n_23), .B(n_24), .ZN(p_1[8]));
   INV_X1 i_34 (.A(p_2[8]), .ZN(n_25));
   OAI22_X1 i_35 (.A1(n_23), .A2(n_24), .B1(n_25), .B2(p_0[8]), .ZN(n_26));
   XNOR2_X1 i_36 (.A(p_0[9]), .B(p_2[9]), .ZN(n_27));
   XNOR2_X1 i_37 (.A(n_26), .B(n_27), .ZN(p_1[9]));
   INV_X1 i_38 (.A(p_0[9]), .ZN(n_28));
   AOI22_X1 i_39 (.A1(n_26), .A2(n_27), .B1(n_28), .B2(p_2[9]), .ZN(n_29));
   XOR2_X1 i_40 (.A(p_0[10]), .B(p_2[10]), .Z(n_30));
   XNOR2_X1 i_41 (.A(n_29), .B(n_30), .ZN(p_1[10]));
   INV_X1 i_42 (.A(p_2[10]), .ZN(n_31));
   OAI22_X1 i_43 (.A1(n_29), .A2(n_30), .B1(n_31), .B2(p_0[10]), .ZN(n_32));
   XNOR2_X1 i_44 (.A(p_0[11]), .B(p_2[11]), .ZN(n_33));
   XNOR2_X1 i_45 (.A(n_32), .B(n_33), .ZN(p_1[11]));
   INV_X1 i_46 (.A(p_0[11]), .ZN(n_34));
   AOI22_X1 i_47 (.A1(n_32), .A2(n_33), .B1(n_34), .B2(p_2[11]), .ZN(n_35));
   XOR2_X1 i_48 (.A(p_0[12]), .B(p_2[12]), .Z(n_36));
   XNOR2_X1 i_49 (.A(n_35), .B(n_36), .ZN(p_1[12]));
   INV_X1 i_50 (.A(p_2[12]), .ZN(n_37));
   OAI22_X1 i_51 (.A1(n_35), .A2(n_36), .B1(n_37), .B2(p_0[12]), .ZN(n_38));
   XNOR2_X1 i_52 (.A(p_0[13]), .B(p_2[13]), .ZN(n_39));
   XNOR2_X1 i_53 (.A(n_38), .B(n_39), .ZN(p_1[13]));
   INV_X1 i_54 (.A(p_0[13]), .ZN(n_40));
   AOI22_X1 i_55 (.A1(n_38), .A2(n_39), .B1(n_40), .B2(p_2[13]), .ZN(n_41));
   INV_X1 i_56 (.A(n_41), .ZN(n_42));
   INV_X1 i_57 (.A(p_2[14]), .ZN(n_43));
   NAND2_X1 i_58 (.A1(n_43), .A2(p_0[14]), .ZN(n_44));
   INV_X1 i_59 (.A(n_44), .ZN(n_45));
   OR2_X1 i_60 (.A1(n_43), .A2(p_0[14]), .ZN(n_46));
   AOI21_X1 i_61 (.A(n_45), .B1(n_41), .B2(n_46), .ZN(n_47));
   NAND2_X1 i_62 (.A1(n_47), .A2(n_46), .ZN(n_48));
   INV_X1 i_63 (.A(n_47), .ZN(n_49));
   AOI22_X1 i_64 (.A1(n_42), .A2(n_48), .B1(n_49), .B2(n_44), .ZN(p_1[14]));
   XNOR2_X1 i_65 (.A(p_0[15]), .B(p_2[15]), .ZN(n_50));
   XNOR2_X1 i_66 (.A(n_47), .B(n_50), .ZN(p_1[15]));
   INV_X1 i_67 (.A(p_0[15]), .ZN(n_51));
   AOI22_X1 i_68 (.A1(n_47), .A2(n_50), .B1(n_51), .B2(p_2[15]), .ZN(n_52));
   XOR2_X1 i_69 (.A(p_0[16]), .B(p_2[16]), .Z(n_53));
   XNOR2_X1 i_70 (.A(n_52), .B(n_53), .ZN(p_1[16]));
   INV_X1 i_71 (.A(p_2[16]), .ZN(n_54));
   OAI22_X1 i_72 (.A1(n_52), .A2(n_53), .B1(n_54), .B2(p_0[16]), .ZN(n_55));
   XNOR2_X1 i_73 (.A(p_0[17]), .B(p_2[17]), .ZN(n_56));
   XNOR2_X1 i_74 (.A(n_55), .B(n_56), .ZN(p_1[17]));
   INV_X1 i_75 (.A(p_0[17]), .ZN(n_57));
   AOI22_X1 i_76 (.A1(n_55), .A2(n_56), .B1(n_57), .B2(p_2[17]), .ZN(n_58));
   XOR2_X1 i_77 (.A(p_0[18]), .B(p_2[18]), .Z(n_59));
   XNOR2_X1 i_78 (.A(n_58), .B(n_59), .ZN(p_1[18]));
   INV_X1 i_79 (.A(p_2[18]), .ZN(n_60));
   OAI22_X1 i_80 (.A1(n_58), .A2(n_59), .B1(n_60), .B2(p_0[18]), .ZN(n_61));
   XNOR2_X1 i_81 (.A(p_0[19]), .B(p_2[19]), .ZN(n_62));
   XNOR2_X1 i_82 (.A(n_61), .B(n_62), .ZN(p_1[19]));
   INV_X1 i_83 (.A(p_0[19]), .ZN(n_63));
   AOI22_X1 i_84 (.A1(n_61), .A2(n_62), .B1(n_63), .B2(p_2[19]), .ZN(n_64));
   INV_X1 i_85 (.A(n_64), .ZN(n_65));
   INV_X1 i_86 (.A(p_2[20]), .ZN(n_66));
   NAND2_X1 i_87 (.A1(n_66), .A2(p_0[20]), .ZN(n_67));
   INV_X1 i_88 (.A(n_67), .ZN(n_68));
   OR2_X1 i_89 (.A1(n_66), .A2(p_0[20]), .ZN(n_69));
   AOI21_X1 i_90 (.A(n_68), .B1(n_64), .B2(n_69), .ZN(n_70));
   NAND2_X1 i_91 (.A1(n_70), .A2(n_69), .ZN(n_71));
   INV_X1 i_92 (.A(n_70), .ZN(n_72));
   AOI22_X1 i_93 (.A1(n_65), .A2(n_71), .B1(n_72), .B2(n_67), .ZN(p_1[20]));
   XNOR2_X1 i_94 (.A(p_0[21]), .B(p_2[21]), .ZN(n_73));
   XNOR2_X1 i_95 (.A(n_70), .B(n_73), .ZN(p_1[21]));
   INV_X1 i_96 (.A(p_0[21]), .ZN(n_74));
   AOI22_X1 i_97 (.A1(n_70), .A2(n_73), .B1(n_74), .B2(p_2[21]), .ZN(n_75));
   XOR2_X1 i_98 (.A(p_0[22]), .B(p_2[22]), .Z(n_76));
   XNOR2_X1 i_99 (.A(n_75), .B(n_76), .ZN(p_1[22]));
   INV_X1 i_100 (.A(p_2[22]), .ZN(n_77));
   OAI22_X1 i_101 (.A1(n_75), .A2(n_76), .B1(n_77), .B2(p_0[22]), .ZN(n_78));
   XOR2_X1 i_102 (.A(p_2[23]), .B(p_0[23]), .Z(n_79));
   XOR2_X1 i_103 (.A(n_78), .B(n_79), .Z(p_1[23]));
   INV_X1 i_104 (.A(n_78), .ZN(n_80));
   INV_X1 i_105 (.A(p_2[23]), .ZN(n_81));
   OAI22_X1 i_106 (.A1(n_80), .A2(n_79), .B1(n_81), .B2(p_0[23]), .ZN(p_1[24]));
endmodule

module adder(a, b, out);
   input [31:0]a;
   input [31:0]b;
   output [31:0]out;

   wire CSA_COUT;
   wire [23:0]CSA_SUM;
   wire [24:0]o_m;
   wire [7:0]o_e;
   wire n_0_6;
   wire n_0_0;
   wire n_0_7;
   wire n_0_1;
   wire n_0_8;
   wire n_0_2;
   wire n_0_9;
   wire n_0_3;
   wire n_0_10;
   wire n_0_4;
   wire n_0_11;
   wire n_0_5;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_317;
   wire n_0_318;
   wire n_0_319;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_332;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_337;
   wire n_0_338;
   wire n_0_339;
   wire n_0_340;
   wire n_0_341;
   wire n_0_342;
   wire n_0_343;
   wire n_0_344;
   wire n_0_345;
   wire n_0_346;
   wire n_0_347;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_355;
   wire n_0_356;
   wire n_0_357;
   wire n_0_358;
   wire n_0_359;
   wire n_0_360;
   wire n_0_361;
   wire n_0_362;
   wire n_0_363;
   wire n_0_364;
   wire n_0_365;
   wire n_0_366;
   wire n_0_367;
   wire n_0_368;
   wire n_0_369;
   wire n_0_370;
   wire n_0_371;
   wire n_0_372;
   wire n_0_373;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_377;
   wire n_0_378;
   wire n_0_379;
   wire n_0_380;
   wire n_0_381;
   wire n_0_382;
   wire n_0_383;
   wire n_0_384;
   wire n_0_385;
   wire n_0_386;
   wire n_0_387;
   wire n_0_388;
   wire n_0_389;
   wire n_0_390;
   wire n_0_391;
   wire n_0_392;
   wire n_0_393;
   wire n_0_394;
   wire n_0_395;
   wire n_0_396;
   wire n_0_397;
   wire n_0_398;
   wire n_0_399;
   wire n_0_400;
   wire n_0_401;
   wire n_0_402;
   wire n_0_403;
   wire n_0_404;
   wire n_0_405;
   wire n_0_406;
   wire n_0_407;
   wire n_0_408;
   wire n_0_409;
   wire n_0_410;
   wire n_0_411;
   wire n_0_412;
   wire n_0_413;
   wire n_0_414;
   wire n_0_415;
   wire n_0_416;
   wire n_0_417;
   wire n_0_418;
   wire n_0_419;
   wire n_0_420;
   wire n_0_421;
   wire n_0_422;
   wire n_0_423;
   wire n_0_424;
   wire n_0_425;
   wire n_0_426;
   wire n_0_427;
   wire n_0_428;
   wire n_0_429;
   wire n_0_430;
   wire n_0_431;
   wire n_0_432;
   wire n_0_433;
   wire n_0_434;
   wire n_0_435;
   wire n_0_436;
   wire n_0_437;
   wire n_0_438;
   wire n_0_439;
   wire n_0_440;
   wire n_0_441;
   wire n_0_442;
   wire n_0_443;
   wire n_0_444;
   wire n_0_445;
   wire n_0_446;
   wire n_0_447;
   wire n_0_448;
   wire n_0_449;
   wire n_0_450;
   wire n_0_451;
   wire n_0_452;
   wire n_0_453;
   wire n_0_454;
   wire n_0_455;
   wire n_0_456;
   wire n_0_457;
   wire n_0_458;
   wire n_0_459;
   wire n_0_460;
   wire n_0_461;
   wire n_0_462;
   wire n_0_463;
   wire n_0_464;
   wire n_0_465;
   wire n_0_466;
   wire n_0_467;
   wire n_0_468;
   wire n_0_469;
   wire n_0_470;
   wire n_0_471;
   wire n_0_472;
   wire n_0_473;
   wire n_0_474;
   wire n_0_475;
   wire n_0_476;
   wire n_0_477;
   wire n_0_478;
   wire n_0_479;
   wire n_0_480;
   wire n_0_481;
   wire n_0_482;
   wire n_0_483;
   wire n_0_484;
   wire n_0_485;
   wire n_0_486;
   wire n_0_487;
   wire n_0_488;
   wire n_0_489;
   wire n_0_490;
   wire n_0_491;
   wire n_0_492;
   wire n_0_493;
   wire n_0_494;
   wire n_0_495;
   wire n_0_496;
   wire n_0_497;
   wire [24:0]i_m;
   wire [7:0]i_e;
   wire [23:0]CSA_IN2;
   wire [23:0]CSA_IN1;

   CSA c1 (.X(CSA_IN1), .Y(CSA_IN2), .Cin(), .S(CSA_SUM), .Cout(CSA_COUT), .OF());
   addition_normaliser norm1 (.in_e(i_e), .in_m({uc_0, i_m[23], i_m[22], i_m[21], 
      i_m[20], i_m[19], i_m[18], i_m[17], i_m[16], i_m[15], i_m[14], i_m[13], 
      i_m[12], i_m[11], i_m[10], i_m[9], i_m[8], i_m[7], i_m[6], i_m[5], i_m[4], 
      i_m[3], i_m[2], i_m[1], i_m[0]}), .out_e(o_e), .out_m({uc_1, uc_2, o_m[22], 
      o_m[21], o_m[20], o_m[19], o_m[18], o_m[17], o_m[16], o_m[15], o_m[14], 
      o_m[13], o_m[12], o_m[11], o_m[10], o_m[9], o_m[8], o_m[7], o_m[6], o_m[5], 
      o_m[4], o_m[3], o_m[2], o_m[1], uc_3}));
   datapath__0_57 i_11 (.p_0({n_155, b[22], b[21], b[20], b[19], b[18], b[17], 
      b[16], b[15], b[14], b[13], b[12], b[11], b[10], b[9], b[8], b[7], b[6], 
      b[5], b[4], b[3], b[2], b[1], b[0]}), .p_1({n_24, n_23, n_22, n_21, n_20, 
      n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, 
      n_6, n_5, n_4, n_3, n_2, n_1, n_0}), .p_2({n_179, n_178, n_177, n_176, 
      n_175, n_174, n_173, n_172, n_171, n_170, n_169, n_168, n_167, n_166, 
      n_165, n_164, n_163, n_162, n_161, n_160, n_159, n_158, n_157, n_156}));
   datapath__0_62 i_16 (.p_0({n_180, a[22], a[21], a[20], a[19], a[18], a[17], 
      a[16], a[15], a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7], a[6], 
      a[5], a[4], a[3], a[2], a[1], a[0]}), .p_1({n_49, n_48, n_47, n_46, n_45, 
      n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, 
      n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25}), .p_2({n_154, n_153, 
      n_152, n_151, n_150, n_149, n_148, n_147, n_146, n_145, n_144, n_143, 
      n_142, n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, n_133, 
      n_132, n_131}));
   HA_X1 i_0_0 (.A(n_124), .B(n_123), .CO(n_0_0), .S(n_0_6));
   HA_X1 i_0_1 (.A(n_125), .B(n_0_0), .CO(n_0_1), .S(n_0_7));
   HA_X1 i_0_2 (.A(n_126), .B(n_0_1), .CO(n_0_2), .S(n_0_8));
   HA_X1 i_0_3 (.A(n_127), .B(n_0_2), .CO(n_0_3), .S(n_0_9));
   HA_X1 i_0_4 (.A(n_128), .B(n_0_3), .CO(n_0_4), .S(n_0_10));
   HA_X1 i_0_5 (.A(n_129), .B(n_0_4), .CO(n_0_5), .S(n_0_11));
   INV_X1 i_0_6 (.A(n_0_12), .ZN(n_50));
   AOI22_X1 i_0_7 (.A1(b[0]), .A2(n_0_187), .B1(a[0]), .B2(n_0_188), .ZN(n_0_12));
   INV_X1 i_0_8 (.A(n_0_13), .ZN(n_51));
   AOI22_X1 i_0_9 (.A1(b[1]), .A2(n_0_187), .B1(a[1]), .B2(n_0_188), .ZN(n_0_13));
   INV_X1 i_0_10 (.A(n_0_14), .ZN(n_52));
   AOI22_X1 i_0_11 (.A1(b[2]), .A2(n_0_187), .B1(a[2]), .B2(n_0_188), .ZN(n_0_14));
   INV_X1 i_0_12 (.A(n_0_15), .ZN(n_53));
   AOI22_X1 i_0_13 (.A1(b[3]), .A2(n_0_187), .B1(a[3]), .B2(n_0_188), .ZN(n_0_15));
   INV_X1 i_0_14 (.A(n_0_16), .ZN(n_54));
   AOI22_X1 i_0_15 (.A1(b[4]), .A2(n_0_187), .B1(a[4]), .B2(n_0_188), .ZN(n_0_16));
   INV_X1 i_0_16 (.A(n_0_17), .ZN(n_55));
   AOI22_X1 i_0_17 (.A1(b[5]), .A2(n_0_187), .B1(a[5]), .B2(n_0_188), .ZN(n_0_17));
   INV_X1 i_0_18 (.A(n_0_18), .ZN(n_56));
   AOI22_X1 i_0_19 (.A1(b[6]), .A2(n_0_187), .B1(a[6]), .B2(n_0_188), .ZN(n_0_18));
   INV_X1 i_0_20 (.A(n_0_19), .ZN(n_57));
   AOI22_X1 i_0_21 (.A1(b[7]), .A2(n_0_187), .B1(a[7]), .B2(n_0_188), .ZN(n_0_19));
   INV_X1 i_0_22 (.A(n_0_20), .ZN(n_58));
   AOI22_X1 i_0_23 (.A1(b[8]), .A2(n_0_187), .B1(a[8]), .B2(n_0_188), .ZN(n_0_20));
   INV_X1 i_0_24 (.A(n_0_21), .ZN(n_59));
   AOI22_X1 i_0_25 (.A1(b[9]), .A2(n_0_187), .B1(a[9]), .B2(n_0_188), .ZN(n_0_21));
   INV_X1 i_0_26 (.A(n_0_22), .ZN(n_60));
   AOI22_X1 i_0_27 (.A1(b[10]), .A2(n_0_187), .B1(a[10]), .B2(n_0_188), .ZN(
      n_0_22));
   INV_X1 i_0_28 (.A(n_0_23), .ZN(n_61));
   AOI22_X1 i_0_29 (.A1(b[11]), .A2(n_0_187), .B1(a[11]), .B2(n_0_188), .ZN(
      n_0_23));
   INV_X1 i_0_30 (.A(n_0_24), .ZN(n_62));
   AOI22_X1 i_0_31 (.A1(b[12]), .A2(n_0_187), .B1(a[12]), .B2(n_0_188), .ZN(
      n_0_24));
   INV_X1 i_0_32 (.A(n_0_25), .ZN(n_63));
   AOI22_X1 i_0_33 (.A1(b[13]), .A2(n_0_187), .B1(a[13]), .B2(n_0_188), .ZN(
      n_0_25));
   INV_X1 i_0_34 (.A(n_0_26), .ZN(n_64));
   AOI22_X1 i_0_35 (.A1(b[14]), .A2(n_0_187), .B1(a[14]), .B2(n_0_188), .ZN(
      n_0_26));
   INV_X1 i_0_36 (.A(n_0_27), .ZN(n_65));
   AOI22_X1 i_0_37 (.A1(b[15]), .A2(n_0_187), .B1(a[15]), .B2(n_0_188), .ZN(
      n_0_27));
   INV_X1 i_0_38 (.A(n_0_28), .ZN(n_66));
   AOI22_X1 i_0_39 (.A1(b[16]), .A2(n_0_187), .B1(a[16]), .B2(n_0_188), .ZN(
      n_0_28));
   INV_X1 i_0_40 (.A(n_0_29), .ZN(n_67));
   AOI22_X1 i_0_41 (.A1(b[17]), .A2(n_0_187), .B1(a[17]), .B2(n_0_188), .ZN(
      n_0_29));
   INV_X1 i_0_42 (.A(n_0_30), .ZN(n_68));
   AOI22_X1 i_0_43 (.A1(b[18]), .A2(n_0_187), .B1(a[18]), .B2(n_0_188), .ZN(
      n_0_30));
   INV_X1 i_0_44 (.A(n_0_31), .ZN(n_69));
   AOI22_X1 i_0_45 (.A1(b[19]), .A2(n_0_187), .B1(a[19]), .B2(n_0_188), .ZN(
      n_0_31));
   INV_X1 i_0_46 (.A(n_0_32), .ZN(n_70));
   AOI22_X1 i_0_47 (.A1(b[20]), .A2(n_0_187), .B1(a[20]), .B2(n_0_188), .ZN(
      n_0_32));
   INV_X1 i_0_48 (.A(n_0_33), .ZN(n_71));
   AOI22_X1 i_0_49 (.A1(b[21]), .A2(n_0_187), .B1(a[21]), .B2(n_0_188), .ZN(
      n_0_33));
   OAI21_X1 i_0_50 (.A(n_0_34), .B1(n_0_481), .B2(n_0_187), .ZN(n_72));
   NAND2_X1 i_0_51 (.A1(b[22]), .A2(n_0_187), .ZN(n_0_34));
   NAND2_X1 i_0_52 (.A1(n_0_477), .A2(n_0_188), .ZN(n_73));
   OAI21_X1 i_0_53 (.A(n_0_35), .B1(n_0_194), .B2(n_0_189), .ZN(n_74));
   AOI22_X1 i_0_54 (.A1(n_156), .A2(n_0_187), .B1(b[0]), .B2(n_0_420), .ZN(
      n_0_35));
   OAI21_X1 i_0_55 (.A(n_0_36), .B1(n_0_199), .B2(n_0_189), .ZN(n_75));
   AOI22_X1 i_0_56 (.A1(n_157), .A2(n_0_187), .B1(b[1]), .B2(n_0_420), .ZN(
      n_0_36));
   OAI21_X1 i_0_57 (.A(n_0_37), .B1(n_0_204), .B2(n_0_189), .ZN(n_76));
   AOI22_X1 i_0_58 (.A1(n_158), .A2(n_0_187), .B1(b[2]), .B2(n_0_420), .ZN(
      n_0_37));
   OAI21_X1 i_0_59 (.A(n_0_38), .B1(n_0_210), .B2(n_0_189), .ZN(n_77));
   AOI22_X1 i_0_60 (.A1(n_159), .A2(n_0_187), .B1(b[3]), .B2(n_0_420), .ZN(
      n_0_38));
   OAI21_X1 i_0_61 (.A(n_0_39), .B1(n_0_215), .B2(n_0_189), .ZN(n_78));
   AOI22_X1 i_0_62 (.A1(n_160), .A2(n_0_187), .B1(b[4]), .B2(n_0_420), .ZN(
      n_0_39));
   OAI21_X1 i_0_63 (.A(n_0_40), .B1(n_0_345), .B2(n_0_188), .ZN(n_79));
   AOI22_X1 i_0_64 (.A1(n_136), .A2(n_0_190), .B1(b[5]), .B2(n_0_420), .ZN(
      n_0_40));
   OAI21_X1 i_0_65 (.A(n_0_41), .B1(n_0_350), .B2(n_0_188), .ZN(n_80));
   AOI22_X1 i_0_66 (.A1(n_137), .A2(n_0_190), .B1(b[6]), .B2(n_0_420), .ZN(
      n_0_41));
   OAI21_X1 i_0_67 (.A(n_0_42), .B1(n_0_356), .B2(n_0_188), .ZN(n_81));
   AOI22_X1 i_0_68 (.A1(b[7]), .A2(n_0_420), .B1(n_138), .B2(n_0_190), .ZN(
      n_0_42));
   OAI21_X1 i_0_69 (.A(n_0_43), .B1(n_0_362), .B2(n_0_188), .ZN(n_82));
   AOI22_X1 i_0_70 (.A1(b[8]), .A2(n_0_420), .B1(n_139), .B2(n_0_190), .ZN(
      n_0_43));
   OAI21_X1 i_0_71 (.A(n_0_44), .B1(n_0_368), .B2(n_0_188), .ZN(n_83));
   AOI22_X1 i_0_72 (.A1(b[9]), .A2(n_0_420), .B1(n_140), .B2(n_0_190), .ZN(
      n_0_44));
   OAI21_X1 i_0_73 (.A(n_0_45), .B1(n_0_373), .B2(n_0_188), .ZN(n_84));
   AOI22_X1 i_0_74 (.A1(b[10]), .A2(n_0_420), .B1(n_141), .B2(n_0_190), .ZN(
      n_0_45));
   OAI21_X1 i_0_75 (.A(n_0_46), .B1(n_0_251), .B2(n_0_189), .ZN(n_85));
   AOI22_X1 i_0_76 (.A1(n_167), .A2(n_0_187), .B1(b[11]), .B2(n_0_420), .ZN(
      n_0_46));
   OAI21_X1 i_0_77 (.A(n_0_47), .B1(n_0_257), .B2(n_0_189), .ZN(n_86));
   AOI22_X1 i_0_78 (.A1(n_168), .A2(n_0_187), .B1(b[12]), .B2(n_0_420), .ZN(
      n_0_47));
   OAI21_X1 i_0_79 (.A(n_0_48), .B1(n_0_260), .B2(n_0_189), .ZN(n_87));
   AOI22_X1 i_0_80 (.A1(n_169), .A2(n_0_187), .B1(b[13]), .B2(n_0_420), .ZN(
      n_0_48));
   OAI21_X1 i_0_81 (.A(n_0_49), .B1(n_0_263), .B2(n_0_189), .ZN(n_88));
   AOI22_X1 i_0_82 (.A1(b[14]), .A2(n_0_420), .B1(n_170), .B2(n_0_187), .ZN(
      n_0_49));
   OAI21_X1 i_0_83 (.A(n_0_50), .B1(n_0_268), .B2(n_0_189), .ZN(n_89));
   AOI22_X1 i_0_84 (.A1(b[15]), .A2(n_0_420), .B1(n_171), .B2(n_0_187), .ZN(
      n_0_50));
   INV_X1 i_0_85 (.A(n_0_51), .ZN(n_90));
   AOI222_X1 i_0_86 (.A1(b[16]), .A2(n_0_420), .B1(n_147), .B2(n_0_190), 
      .C1(n_172), .C2(n_0_187), .ZN(n_0_51));
   OAI21_X1 i_0_87 (.A(n_0_52), .B1(n_0_278), .B2(n_0_189), .ZN(n_91));
   AOI22_X1 i_0_88 (.A1(n_173), .A2(n_0_187), .B1(b[17]), .B2(n_0_420), .ZN(
      n_0_52));
   OAI21_X1 i_0_89 (.A(n_0_53), .B1(n_0_281), .B2(n_0_189), .ZN(n_92));
   AOI22_X1 i_0_90 (.A1(b[18]), .A2(n_0_420), .B1(n_174), .B2(n_0_187), .ZN(
      n_0_53));
   OAI21_X1 i_0_91 (.A(n_0_54), .B1(n_0_284), .B2(n_0_189), .ZN(n_93));
   AOI22_X1 i_0_92 (.A1(b[19]), .A2(n_0_420), .B1(n_175), .B2(n_0_187), .ZN(
      n_0_54));
   INV_X1 i_0_93 (.A(n_0_55), .ZN(n_94));
   AOI222_X1 i_0_94 (.A1(b[20]), .A2(n_0_420), .B1(n_151), .B2(n_0_190), 
      .C1(n_176), .C2(n_0_187), .ZN(n_0_55));
   INV_X1 i_0_95 (.A(n_0_56), .ZN(n_95));
   AOI222_X1 i_0_96 (.A1(b[21]), .A2(n_0_420), .B1(n_152), .B2(n_0_190), 
      .C1(n_177), .C2(n_0_187), .ZN(n_0_56));
   NAND2_X1 i_0_97 (.A1(n_0_415), .A2(n_0_300), .ZN(n_96));
   INV_X1 i_0_98 (.A(n_0_57), .ZN(n_97));
   AOI222_X1 i_0_99 (.A1(n_25), .A2(n_0_168), .B1(n_0), .B2(n_0_182), .C1(
      CSA_SUM[0]), .C2(n_122), .ZN(n_0_57));
   INV_X1 i_0_100 (.A(n_0_58), .ZN(n_98));
   AOI221_X1 i_0_101 (.A(n_0_86), .B1(n_26), .B2(n_0_168), .C1(CSA_SUM[1]), 
      .C2(n_122), .ZN(n_0_58));
   INV_X1 i_0_102 (.A(n_0_59), .ZN(n_99));
   AOI222_X1 i_0_103 (.A1(n_27), .A2(n_0_168), .B1(CSA_SUM[2]), .B2(n_122), 
      .C1(n_2), .C2(n_0_182), .ZN(n_0_59));
   INV_X1 i_0_104 (.A(n_0_60), .ZN(n_100));
   AOI222_X1 i_0_105 (.A1(n_28), .A2(n_0_168), .B1(CSA_SUM[3]), .B2(n_122), 
      .C1(n_3), .C2(n_0_182), .ZN(n_0_60));
   INV_X1 i_0_106 (.A(n_0_61), .ZN(n_101));
   AOI222_X1 i_0_107 (.A1(n_29), .A2(n_0_168), .B1(CSA_SUM[4]), .B2(n_122), 
      .C1(n_4), .C2(n_0_182), .ZN(n_0_61));
   INV_X1 i_0_108 (.A(n_0_62), .ZN(n_102));
   AOI222_X1 i_0_109 (.A1(n_30), .A2(n_0_168), .B1(CSA_SUM[5]), .B2(n_122), 
      .C1(n_5), .C2(n_0_182), .ZN(n_0_62));
   INV_X1 i_0_110 (.A(n_0_63), .ZN(n_103));
   AOI222_X1 i_0_111 (.A1(n_31), .A2(n_0_168), .B1(CSA_SUM[6]), .B2(n_122), 
      .C1(n_6), .C2(n_0_182), .ZN(n_0_63));
   INV_X1 i_0_112 (.A(n_0_64), .ZN(n_104));
   AOI222_X1 i_0_113 (.A1(n_32), .A2(n_0_168), .B1(CSA_SUM[7]), .B2(n_122), 
      .C1(n_7), .C2(n_0_182), .ZN(n_0_64));
   INV_X1 i_0_114 (.A(n_0_65), .ZN(n_105));
   AOI222_X1 i_0_115 (.A1(n_33), .A2(n_0_168), .B1(CSA_SUM[8]), .B2(n_122), 
      .C1(n_8), .C2(n_0_182), .ZN(n_0_65));
   INV_X1 i_0_116 (.A(n_0_66), .ZN(n_106));
   AOI222_X1 i_0_117 (.A1(n_34), .A2(n_0_168), .B1(CSA_SUM[9]), .B2(n_122), 
      .C1(n_9), .C2(n_0_182), .ZN(n_0_66));
   INV_X1 i_0_118 (.A(n_0_67), .ZN(n_107));
   AOI222_X1 i_0_119 (.A1(n_35), .A2(n_0_168), .B1(CSA_SUM[10]), .B2(n_122), 
      .C1(n_10), .C2(n_0_182), .ZN(n_0_67));
   INV_X1 i_0_120 (.A(n_0_68), .ZN(n_108));
   AOI222_X1 i_0_121 (.A1(n_36), .A2(n_0_168), .B1(CSA_SUM[11]), .B2(n_122), 
      .C1(n_11), .C2(n_0_182), .ZN(n_0_68));
   INV_X1 i_0_122 (.A(n_0_69), .ZN(n_109));
   AOI222_X1 i_0_123 (.A1(n_37), .A2(n_0_168), .B1(CSA_SUM[12]), .B2(n_122), 
      .C1(n_12), .C2(n_0_182), .ZN(n_0_69));
   INV_X1 i_0_124 (.A(n_0_70), .ZN(n_110));
   AOI222_X1 i_0_125 (.A1(n_38), .A2(n_0_168), .B1(CSA_SUM[13]), .B2(n_122), 
      .C1(n_13), .C2(n_0_182), .ZN(n_0_70));
   INV_X1 i_0_126 (.A(n_0_71), .ZN(n_111));
   AOI222_X1 i_0_127 (.A1(n_39), .A2(n_0_168), .B1(CSA_SUM[14]), .B2(n_122), 
      .C1(n_14), .C2(n_0_182), .ZN(n_0_71));
   INV_X1 i_0_128 (.A(n_0_72), .ZN(n_112));
   AOI222_X1 i_0_129 (.A1(n_40), .A2(n_0_168), .B1(CSA_SUM[15]), .B2(n_122), 
      .C1(n_15), .C2(n_0_182), .ZN(n_0_72));
   INV_X1 i_0_130 (.A(n_0_73), .ZN(n_113));
   AOI222_X1 i_0_131 (.A1(n_41), .A2(n_0_168), .B1(CSA_SUM[16]), .B2(n_122), 
      .C1(n_16), .C2(n_0_182), .ZN(n_0_73));
   INV_X1 i_0_132 (.A(n_0_74), .ZN(n_114));
   AOI222_X1 i_0_133 (.A1(n_42), .A2(n_0_168), .B1(CSA_SUM[17]), .B2(n_122), 
      .C1(n_17), .C2(n_0_182), .ZN(n_0_74));
   INV_X1 i_0_134 (.A(n_0_75), .ZN(n_115));
   AOI222_X1 i_0_135 (.A1(n_43), .A2(n_0_168), .B1(CSA_SUM[18]), .B2(n_122), 
      .C1(n_18), .C2(n_0_182), .ZN(n_0_75));
   INV_X1 i_0_136 (.A(n_0_76), .ZN(n_116));
   AOI222_X1 i_0_137 (.A1(n_44), .A2(n_0_168), .B1(CSA_SUM[19]), .B2(n_122), 
      .C1(n_19), .C2(n_0_182), .ZN(n_0_76));
   INV_X1 i_0_138 (.A(n_0_77), .ZN(n_117));
   AOI222_X1 i_0_139 (.A1(n_45), .A2(n_0_168), .B1(CSA_SUM[20]), .B2(n_122), 
      .C1(n_20), .C2(n_0_182), .ZN(n_0_77));
   INV_X1 i_0_140 (.A(n_0_78), .ZN(n_118));
   AOI222_X1 i_0_141 (.A1(n_46), .A2(n_0_168), .B1(CSA_SUM[21]), .B2(n_122), 
      .C1(n_21), .C2(n_0_182), .ZN(n_0_78));
   INV_X1 i_0_142 (.A(n_0_79), .ZN(n_119));
   AOI221_X1 i_0_143 (.A(n_0_152), .B1(n_47), .B2(n_0_168), .C1(CSA_SUM[22]), 
      .C2(n_122), .ZN(n_0_79));
   NAND3_X1 i_0_144 (.A1(n_0_82), .A2(n_0_81), .A3(n_0_80), .ZN(out[0]));
   AOI222_X1 i_0_145 (.A1(n_1), .A2(n_0_171), .B1(n_0), .B2(n_0_179), .C1(
      CSA_SUM[0]), .C2(n_0_150), .ZN(n_0_80));
   NAND2_X1 i_0_146 (.A1(n_25), .A2(n_0_148), .ZN(n_0_81));
   AOI22_X1 i_0_147 (.A1(CSA_SUM[1]), .A2(n_0_169), .B1(n_26), .B2(n_0_166), 
      .ZN(n_0_82));
   NAND3_X1 i_0_148 (.A1(n_0_85), .A2(n_0_83), .A3(n_0_84), .ZN(out[1]));
   AOI222_X1 i_0_149 (.A1(o_m[1]), .A2(n_120), .B1(n_26), .B2(n_0_148), .C1(n_2), 
      .C2(n_0_171), .ZN(n_0_83));
   AOI222_X1 i_0_150 (.A1(n_0_153), .A2(n_0_86), .B1(CSA_SUM[1]), .B2(n_0_150), 
      .C1(n_27), .C2(n_0_166), .ZN(n_0_84));
   NAND2_X1 i_0_151 (.A1(CSA_SUM[2]), .A2(n_0_169), .ZN(n_0_85));
   AND2_X1 i_0_152 (.A1(n_1), .A2(n_0_182), .ZN(n_0_86));
   NAND3_X1 i_0_153 (.A1(n_0_88), .A2(n_0_87), .A3(n_0_89), .ZN(out[2]));
   AOI222_X1 i_0_154 (.A1(n_2), .A2(n_0_179), .B1(CSA_SUM[2]), .B2(n_0_150), 
      .C1(n_28), .C2(n_0_166), .ZN(n_0_87));
   AOI22_X1 i_0_155 (.A1(n_27), .A2(n_0_148), .B1(o_m[2]), .B2(n_120), .ZN(
      n_0_88));
   AOI22_X1 i_0_156 (.A1(n_3), .A2(n_0_171), .B1(CSA_SUM[3]), .B2(n_0_169), 
      .ZN(n_0_89));
   NAND3_X1 i_0_157 (.A1(n_0_91), .A2(n_0_90), .A3(n_0_92), .ZN(out[3]));
   AOI222_X1 i_0_158 (.A1(n_3), .A2(n_0_179), .B1(CSA_SUM[3]), .B2(n_0_150), 
      .C1(n_29), .C2(n_0_166), .ZN(n_0_90));
   AOI22_X1 i_0_159 (.A1(n_28), .A2(n_0_148), .B1(o_m[3]), .B2(n_120), .ZN(
      n_0_91));
   AOI22_X1 i_0_160 (.A1(n_4), .A2(n_0_171), .B1(CSA_SUM[4]), .B2(n_0_169), 
      .ZN(n_0_92));
   NAND3_X1 i_0_161 (.A1(n_0_94), .A2(n_0_93), .A3(n_0_95), .ZN(out[4]));
   AOI222_X1 i_0_162 (.A1(n_4), .A2(n_0_179), .B1(CSA_SUM[4]), .B2(n_0_150), 
      .C1(n_30), .C2(n_0_166), .ZN(n_0_93));
   AOI22_X1 i_0_163 (.A1(n_29), .A2(n_0_148), .B1(o_m[4]), .B2(n_120), .ZN(
      n_0_94));
   AOI22_X1 i_0_164 (.A1(n_5), .A2(n_0_171), .B1(CSA_SUM[5]), .B2(n_0_169), 
      .ZN(n_0_95));
   NAND3_X1 i_0_165 (.A1(n_0_97), .A2(n_0_96), .A3(n_0_98), .ZN(out[5]));
   AOI222_X1 i_0_166 (.A1(n_5), .A2(n_0_179), .B1(CSA_SUM[5]), .B2(n_0_150), 
      .C1(n_31), .C2(n_0_166), .ZN(n_0_96));
   AOI22_X1 i_0_167 (.A1(n_30), .A2(n_0_148), .B1(o_m[5]), .B2(n_120), .ZN(
      n_0_97));
   AOI22_X1 i_0_168 (.A1(n_6), .A2(n_0_171), .B1(CSA_SUM[6]), .B2(n_0_169), 
      .ZN(n_0_98));
   NAND3_X1 i_0_169 (.A1(n_0_100), .A2(n_0_99), .A3(n_0_101), .ZN(out[6]));
   AOI222_X1 i_0_170 (.A1(n_6), .A2(n_0_179), .B1(CSA_SUM[6]), .B2(n_0_150), 
      .C1(n_32), .C2(n_0_166), .ZN(n_0_99));
   AOI22_X1 i_0_171 (.A1(n_31), .A2(n_0_148), .B1(o_m[6]), .B2(n_120), .ZN(
      n_0_100));
   AOI22_X1 i_0_172 (.A1(n_7), .A2(n_0_171), .B1(CSA_SUM[7]), .B2(n_0_169), 
      .ZN(n_0_101));
   NAND3_X1 i_0_173 (.A1(n_0_103), .A2(n_0_102), .A3(n_0_104), .ZN(out[7]));
   AOI222_X1 i_0_174 (.A1(n_7), .A2(n_0_179), .B1(CSA_SUM[7]), .B2(n_0_150), 
      .C1(n_33), .C2(n_0_166), .ZN(n_0_102));
   AOI22_X1 i_0_175 (.A1(n_32), .A2(n_0_148), .B1(o_m[7]), .B2(n_120), .ZN(
      n_0_103));
   AOI22_X1 i_0_176 (.A1(n_8), .A2(n_0_171), .B1(CSA_SUM[8]), .B2(n_0_169), 
      .ZN(n_0_104));
   NAND3_X1 i_0_177 (.A1(n_0_106), .A2(n_0_105), .A3(n_0_107), .ZN(out[8]));
   AOI222_X1 i_0_178 (.A1(n_8), .A2(n_0_179), .B1(CSA_SUM[8]), .B2(n_0_150), 
      .C1(n_34), .C2(n_0_166), .ZN(n_0_105));
   AOI22_X1 i_0_179 (.A1(n_33), .A2(n_0_148), .B1(o_m[8]), .B2(n_120), .ZN(
      n_0_106));
   AOI22_X1 i_0_180 (.A1(n_9), .A2(n_0_171), .B1(CSA_SUM[9]), .B2(n_0_169), 
      .ZN(n_0_107));
   NAND3_X1 i_0_181 (.A1(n_0_109), .A2(n_0_108), .A3(n_0_110), .ZN(out[9]));
   AOI222_X1 i_0_182 (.A1(n_9), .A2(n_0_179), .B1(CSA_SUM[9]), .B2(n_0_150), 
      .C1(n_35), .C2(n_0_166), .ZN(n_0_108));
   AOI22_X1 i_0_183 (.A1(n_34), .A2(n_0_148), .B1(o_m[9]), .B2(n_120), .ZN(
      n_0_109));
   AOI22_X1 i_0_184 (.A1(n_10), .A2(n_0_171), .B1(CSA_SUM[10]), .B2(n_0_169), 
      .ZN(n_0_110));
   NAND3_X1 i_0_185 (.A1(n_0_112), .A2(n_0_111), .A3(n_0_113), .ZN(out[10]));
   AOI222_X1 i_0_186 (.A1(n_10), .A2(n_0_179), .B1(CSA_SUM[10]), .B2(n_0_150), 
      .C1(n_36), .C2(n_0_166), .ZN(n_0_111));
   AOI22_X1 i_0_187 (.A1(n_35), .A2(n_0_148), .B1(o_m[10]), .B2(n_120), .ZN(
      n_0_112));
   AOI22_X1 i_0_188 (.A1(n_11), .A2(n_0_171), .B1(CSA_SUM[11]), .B2(n_0_169), 
      .ZN(n_0_113));
   NAND3_X1 i_0_189 (.A1(n_0_115), .A2(n_0_114), .A3(n_0_116), .ZN(out[11]));
   AOI222_X1 i_0_190 (.A1(n_11), .A2(n_0_179), .B1(CSA_SUM[11]), .B2(n_0_150), 
      .C1(n_37), .C2(n_0_166), .ZN(n_0_114));
   AOI22_X1 i_0_191 (.A1(n_36), .A2(n_0_148), .B1(o_m[11]), .B2(n_120), .ZN(
      n_0_115));
   AOI22_X1 i_0_192 (.A1(n_12), .A2(n_0_171), .B1(CSA_SUM[12]), .B2(n_0_169), 
      .ZN(n_0_116));
   NAND3_X1 i_0_193 (.A1(n_0_118), .A2(n_0_117), .A3(n_0_119), .ZN(out[12]));
   AOI222_X1 i_0_194 (.A1(n_12), .A2(n_0_179), .B1(CSA_SUM[12]), .B2(n_0_150), 
      .C1(n_38), .C2(n_0_166), .ZN(n_0_117));
   AOI22_X1 i_0_195 (.A1(n_37), .A2(n_0_148), .B1(o_m[12]), .B2(n_120), .ZN(
      n_0_118));
   AOI22_X1 i_0_196 (.A1(n_13), .A2(n_0_171), .B1(CSA_SUM[13]), .B2(n_0_169), 
      .ZN(n_0_119));
   NAND3_X1 i_0_197 (.A1(n_0_121), .A2(n_0_120), .A3(n_0_122), .ZN(out[13]));
   AOI222_X1 i_0_198 (.A1(n_13), .A2(n_0_179), .B1(CSA_SUM[13]), .B2(n_0_150), 
      .C1(n_39), .C2(n_0_166), .ZN(n_0_120));
   AOI22_X1 i_0_199 (.A1(n_38), .A2(n_0_148), .B1(o_m[13]), .B2(n_120), .ZN(
      n_0_121));
   AOI22_X1 i_0_200 (.A1(n_14), .A2(n_0_171), .B1(CSA_SUM[14]), .B2(n_0_169), 
      .ZN(n_0_122));
   NAND3_X1 i_0_201 (.A1(n_0_124), .A2(n_0_123), .A3(n_0_125), .ZN(out[14]));
   AOI222_X1 i_0_202 (.A1(n_14), .A2(n_0_179), .B1(CSA_SUM[14]), .B2(n_0_150), 
      .C1(n_40), .C2(n_0_166), .ZN(n_0_123));
   AOI22_X1 i_0_203 (.A1(n_39), .A2(n_0_148), .B1(o_m[14]), .B2(n_120), .ZN(
      n_0_124));
   AOI22_X1 i_0_204 (.A1(n_15), .A2(n_0_171), .B1(CSA_SUM[15]), .B2(n_0_169), 
      .ZN(n_0_125));
   NAND3_X1 i_0_205 (.A1(n_0_127), .A2(n_0_126), .A3(n_0_128), .ZN(out[15]));
   AOI222_X1 i_0_206 (.A1(n_15), .A2(n_0_179), .B1(CSA_SUM[15]), .B2(n_0_150), 
      .C1(n_41), .C2(n_0_166), .ZN(n_0_126));
   AOI22_X1 i_0_207 (.A1(n_40), .A2(n_0_148), .B1(o_m[15]), .B2(n_120), .ZN(
      n_0_127));
   AOI22_X1 i_0_208 (.A1(n_16), .A2(n_0_171), .B1(CSA_SUM[16]), .B2(n_0_169), 
      .ZN(n_0_128));
   NAND3_X1 i_0_209 (.A1(n_0_130), .A2(n_0_129), .A3(n_0_131), .ZN(out[16]));
   AOI222_X1 i_0_210 (.A1(n_16), .A2(n_0_179), .B1(CSA_SUM[16]), .B2(n_0_150), 
      .C1(n_42), .C2(n_0_166), .ZN(n_0_129));
   AOI22_X1 i_0_211 (.A1(n_41), .A2(n_0_148), .B1(o_m[16]), .B2(n_120), .ZN(
      n_0_130));
   AOI22_X1 i_0_212 (.A1(n_17), .A2(n_0_171), .B1(CSA_SUM[17]), .B2(n_0_169), 
      .ZN(n_0_131));
   NAND3_X1 i_0_213 (.A1(n_0_133), .A2(n_0_132), .A3(n_0_134), .ZN(out[17]));
   AOI222_X1 i_0_214 (.A1(n_17), .A2(n_0_179), .B1(CSA_SUM[17]), .B2(n_0_150), 
      .C1(n_43), .C2(n_0_166), .ZN(n_0_132));
   AOI22_X1 i_0_215 (.A1(n_42), .A2(n_0_148), .B1(o_m[17]), .B2(n_120), .ZN(
      n_0_133));
   AOI22_X1 i_0_216 (.A1(n_18), .A2(n_0_171), .B1(CSA_SUM[18]), .B2(n_0_169), 
      .ZN(n_0_134));
   NAND3_X1 i_0_217 (.A1(n_0_136), .A2(n_0_135), .A3(n_0_137), .ZN(out[18]));
   AOI222_X1 i_0_218 (.A1(n_18), .A2(n_0_179), .B1(CSA_SUM[18]), .B2(n_0_150), 
      .C1(n_44), .C2(n_0_166), .ZN(n_0_135));
   AOI22_X1 i_0_219 (.A1(n_43), .A2(n_0_148), .B1(o_m[18]), .B2(n_120), .ZN(
      n_0_136));
   AOI22_X1 i_0_220 (.A1(n_19), .A2(n_0_171), .B1(CSA_SUM[19]), .B2(n_0_169), 
      .ZN(n_0_137));
   NAND3_X1 i_0_221 (.A1(n_0_139), .A2(n_0_138), .A3(n_0_140), .ZN(out[19]));
   AOI222_X1 i_0_222 (.A1(n_19), .A2(n_0_179), .B1(CSA_SUM[19]), .B2(n_0_150), 
      .C1(n_45), .C2(n_0_166), .ZN(n_0_138));
   AOI22_X1 i_0_223 (.A1(n_44), .A2(n_0_148), .B1(o_m[19]), .B2(n_120), .ZN(
      n_0_139));
   AOI22_X1 i_0_224 (.A1(n_20), .A2(n_0_171), .B1(CSA_SUM[20]), .B2(n_0_169), 
      .ZN(n_0_140));
   NAND3_X1 i_0_225 (.A1(n_0_142), .A2(n_0_141), .A3(n_0_143), .ZN(out[20]));
   AOI222_X1 i_0_226 (.A1(n_20), .A2(n_0_179), .B1(CSA_SUM[20]), .B2(n_0_150), 
      .C1(n_46), .C2(n_0_166), .ZN(n_0_141));
   AOI22_X1 i_0_227 (.A1(n_45), .A2(n_0_148), .B1(o_m[20]), .B2(n_120), .ZN(
      n_0_142));
   AOI22_X1 i_0_228 (.A1(n_21), .A2(n_0_171), .B1(CSA_SUM[21]), .B2(n_0_169), 
      .ZN(n_0_143));
   NAND3_X1 i_0_229 (.A1(n_0_145), .A2(n_0_144), .A3(n_0_146), .ZN(out[21]));
   AOI222_X1 i_0_230 (.A1(n_21), .A2(n_0_179), .B1(CSA_SUM[21]), .B2(n_0_150), 
      .C1(n_47), .C2(n_0_166), .ZN(n_0_144));
   AOI22_X1 i_0_231 (.A1(n_46), .A2(n_0_148), .B1(o_m[21]), .B2(n_120), .ZN(
      n_0_145));
   AOI22_X1 i_0_232 (.A1(n_22), .A2(n_0_171), .B1(CSA_SUM[22]), .B2(n_0_169), 
      .ZN(n_0_146));
   NAND3_X1 i_0_233 (.A1(n_0_149), .A2(n_0_147), .A3(n_0_151), .ZN(out[22]));
   AOI222_X1 i_0_234 (.A1(o_m[22]), .A2(n_120), .B1(n_47), .B2(n_0_148), 
      .C1(n_48), .C2(n_0_166), .ZN(n_0_147));
   AND2_X1 i_0_235 (.A1(n_0_168), .A2(n_0_153), .ZN(n_0_148));
   AOI22_X1 i_0_236 (.A1(n_0_153), .A2(n_0_152), .B1(CSA_SUM[22]), .B2(n_0_150), 
      .ZN(n_0_149));
   AND2_X1 i_0_237 (.A1(n_0_184), .A2(n_0_153), .ZN(n_0_150));
   AOI22_X1 i_0_238 (.A1(n_24), .A2(n_0_180), .B1(CSA_SUM[23]), .B2(n_0_169), 
      .ZN(n_0_151));
   AND2_X1 i_0_239 (.A1(n_22), .A2(n_0_182), .ZN(n_0_152));
   NOR2_X1 i_0_240 (.A1(n_0_165), .A2(n_0_163), .ZN(n_0_153));
   OAI221_X1 i_0_241 (.A(n_0_154), .B1(n_123), .B2(n_0_164), .C1(n_0_473), 
      .C2(n_0_177), .ZN(out[23]));
   AOI22_X1 i_0_242 (.A1(o_e[0]), .A2(n_120), .B1(n_0_472), .B2(n_0_173), 
      .ZN(n_0_154));
   OAI21_X1 i_0_243 (.A(n_0_155), .B1(n_0_490), .B2(n_0_177), .ZN(out[24]));
   AOI222_X1 i_0_244 (.A1(o_e[1]), .A2(n_120), .B1(n_0_6), .B2(n_0_165), 
      .C1(a[24]), .C2(n_0_173), .ZN(n_0_155));
   OAI21_X1 i_0_245 (.A(n_0_156), .B1(n_0_491), .B2(n_0_177), .ZN(out[25]));
   AOI222_X1 i_0_246 (.A1(o_e[2]), .A2(n_120), .B1(n_0_7), .B2(n_0_165), 
      .C1(a[25]), .C2(n_0_173), .ZN(n_0_156));
   OAI21_X1 i_0_247 (.A(n_0_157), .B1(n_0_492), .B2(n_0_177), .ZN(out[26]));
   AOI222_X1 i_0_248 (.A1(o_e[3]), .A2(n_120), .B1(n_0_8), .B2(n_0_165), 
      .C1(a[26]), .C2(n_0_173), .ZN(n_0_157));
   OAI21_X1 i_0_249 (.A(n_0_158), .B1(n_0_493), .B2(n_0_177), .ZN(out[27]));
   AOI222_X1 i_0_250 (.A1(o_e[4]), .A2(n_120), .B1(n_0_9), .B2(n_0_165), 
      .C1(a[27]), .C2(n_0_173), .ZN(n_0_158));
   OAI21_X1 i_0_251 (.A(n_0_159), .B1(n_0_494), .B2(n_0_177), .ZN(out[28]));
   AOI222_X1 i_0_252 (.A1(o_e[5]), .A2(n_120), .B1(n_0_10), .B2(n_0_165), 
      .C1(a[28]), .C2(n_0_173), .ZN(n_0_159));
   OAI21_X1 i_0_253 (.A(n_0_160), .B1(n_0_495), .B2(n_0_177), .ZN(out[29]));
   AOI222_X1 i_0_254 (.A1(o_e[6]), .A2(n_120), .B1(n_0_11), .B2(n_0_165), 
      .C1(a[29]), .C2(n_0_173), .ZN(n_0_160));
   OAI21_X1 i_0_255 (.A(n_0_161), .B1(n_0_496), .B2(n_0_177), .ZN(out[30]));
   AOI221_X1 i_0_256 (.A(n_0_162), .B1(o_e[7]), .B2(n_120), .C1(a[30]), .C2(
      n_0_173), .ZN(n_0_161));
   AOI221_X1 i_0_257 (.A(n_0_164), .B1(n_0_480), .B2(n_0_193), .C1(n_0_5), 
      .C2(n_130), .ZN(n_0_162));
   NOR2_X1 i_0_258 (.A1(n_0_165), .A2(n_121), .ZN(n_120));
   INV_X1 i_0_259 (.A(n_0_163), .ZN(n_121));
   AOI221_X1 i_0_260 (.A(n_0_180), .B1(CSA_SUM[23]), .B2(n_122), .C1(n_48), 
      .C2(n_0_168), .ZN(n_0_163));
   INV_X1 i_0_261 (.A(n_0_165), .ZN(n_0_164));
   NAND3_X1 i_0_262 (.A1(n_0_170), .A2(n_0_167), .A3(n_0_172), .ZN(n_0_165));
   INV_X1 i_0_263 (.A(n_0_167), .ZN(n_0_166));
   NAND2_X1 i_0_264 (.A1(n_49), .A2(n_0_168), .ZN(n_0_167));
   NOR2_X1 i_0_265 (.A1(n_0_189), .A2(n_0_184), .ZN(n_0_168));
   INV_X1 i_0_266 (.A(n_0_170), .ZN(n_0_169));
   AOI21_X1 i_0_267 (.A(n_0_420), .B1(CSA_COUT), .B2(n_0_184), .ZN(n_0_170));
   INV_X1 i_0_268 (.A(n_0_172), .ZN(n_0_171));
   NAND2_X1 i_0_269 (.A1(n_24), .A2(n_0_182), .ZN(n_0_172));
   AOI211_X1 i_0_270 (.A(n_0_174), .B(n_0_176), .C1(n_49), .C2(n_0_183), 
      .ZN(n_0_173));
   INV_X1 i_0_271 (.A(n_0_175), .ZN(n_0_174));
   AOI21_X1 i_0_272 (.A(n_0_189), .B1(CSA_COUT), .B2(n_0_184), .ZN(n_0_175));
   AOI221_X1 i_0_273 (.A(n_0_420), .B1(n_48), .B2(n_0_183), .C1(CSA_SUM[23]), 
      .C2(n_0_184), .ZN(n_0_176));
   AOI21_X1 i_0_274 (.A(n_0_179), .B1(CSA_SUM[23]), .B2(n_0_178), .ZN(n_0_177));
   NOR3_X1 i_0_275 (.A1(CSA_COUT), .A2(n_0_183), .A3(n_0_188), .ZN(n_0_178));
   NOR2_X1 i_0_276 (.A1(n_24), .A2(n_0_181), .ZN(n_0_179));
   INV_X1 i_0_277 (.A(n_0_181), .ZN(n_0_180));
   NAND2_X1 i_0_278 (.A1(n_23), .A2(n_0_182), .ZN(n_0_181));
   NOR2_X1 i_0_279 (.A1(n_0_190), .A2(n_122), .ZN(n_0_182));
   NAND2_X1 i_0_280 (.A1(n_0_421), .A2(n_0_183), .ZN(n_122));
   INV_X1 i_0_281 (.A(n_0_184), .ZN(n_0_183));
   AOI22_X1 i_0_282 (.A1(n_0_497), .A2(a[31]), .B1(b[31]), .B2(n_0_488), 
      .ZN(n_0_184));
   OAI22_X1 i_0_283 (.A1(n_0_497), .A2(n_0_188), .B1(n_0_488), .B2(n_0_187), 
      .ZN(out[31]));
   AOI22_X1 i_0_284 (.A1(n_0_473), .A2(n_0_189), .B1(n_0_471), .B2(n_0_190), 
      .ZN(n_123));
   OAI21_X1 i_0_285 (.A(n_0_185), .B1(n_0_490), .B2(n_0_188), .ZN(n_124));
   NAND2_X1 i_0_286 (.A1(a[24]), .A2(n_0_188), .ZN(n_0_185));
   OAI22_X1 i_0_287 (.A1(n_0_491), .A2(n_0_188), .B1(n_0_483), .B2(n_0_187), 
      .ZN(n_125));
   OAI22_X1 i_0_288 (.A1(n_0_492), .A2(n_0_188), .B1(n_0_484), .B2(n_0_187), 
      .ZN(n_126));
   OAI21_X1 i_0_289 (.A(n_0_186), .B1(n_0_493), .B2(n_0_188), .ZN(n_127));
   NAND2_X1 i_0_290 (.A1(a[27]), .A2(n_0_188), .ZN(n_0_186));
   OAI22_X1 i_0_291 (.A1(n_0_494), .A2(n_0_188), .B1(n_0_485), .B2(n_0_187), 
      .ZN(n_128));
   OAI22_X1 i_0_292 (.A1(n_0_495), .A2(n_0_188), .B1(n_0_486), .B2(n_0_187), 
      .ZN(n_129));
   INV_X1 i_0_293 (.A(n_0_188), .ZN(n_0_187));
   NAND2_X1 i_0_294 (.A1(n_0_421), .A2(n_0_189), .ZN(n_0_188));
   INV_X1 i_0_295 (.A(n_0_190), .ZN(n_0_189));
   AOI22_X1 i_0_296 (.A1(b[30]), .A2(n_0_487), .B1(n_0_445), .B2(n_0_191), 
      .ZN(n_0_190));
   AOI22_X1 i_0_297 (.A1(n_0_496), .A2(a[30]), .B1(n_0_446), .B2(n_0_192), 
      .ZN(n_0_191));
   AOI21_X1 i_0_298 (.A(n_0_447), .B1(n_0_449), .B2(n_0_440), .ZN(n_0_192));
   INV_X1 i_0_299 (.A(n_130), .ZN(n_0_193));
   NAND2_X1 i_0_300 (.A1(n_0_496), .A2(n_0_487), .ZN(n_130));
   INV_X1 i_0_301 (.A(n_0_194), .ZN(n_131));
   AOI22_X1 i_0_302 (.A1(n_0_286), .A2(n_0_200), .B1(n_0_287), .B2(n_0_195), 
      .ZN(n_0_194));
   AOI22_X1 i_0_303 (.A1(n_0_303), .A2(n_0_206), .B1(n_0_302), .B2(n_0_196), 
      .ZN(n_0_195));
   AOI221_X1 i_0_304 (.A(n_0_197), .B1(b[0]), .B2(n_0_305), .C1(n_0_306), 
      .C2(n_0_218), .ZN(n_0_196));
   NOR2_X1 i_0_305 (.A1(n_0_306), .A2(n_0_198), .ZN(n_0_197));
   AOI22_X1 i_0_306 (.A1(b[16]), .A2(n_0_235), .B1(b[8]), .B2(n_0_274), .ZN(
      n_0_198));
   INV_X1 i_0_307 (.A(n_0_199), .ZN(n_132));
   AOI22_X1 i_0_308 (.A1(n_0_286), .A2(n_0_205), .B1(n_0_287), .B2(n_0_200), 
      .ZN(n_0_199));
   INV_X1 i_0_309 (.A(n_0_201), .ZN(n_0_200));
   AOI21_X1 i_0_310 (.A(n_0_202), .B1(n_0_303), .B2(n_0_213), .ZN(n_0_201));
   AOI221_X1 i_0_311 (.A(n_0_303), .B1(n_0_307), .B2(n_0_203), .C1(n_0_306), 
      .C2(n_0_224), .ZN(n_0_202));
   AOI222_X1 i_0_312 (.A1(b[1]), .A2(n_0_308), .B1(b[9]), .B2(n_0_274), .C1(
      b[17]), .C2(n_0_235), .ZN(n_0_203));
   INV_X1 i_0_313 (.A(n_0_204), .ZN(n_133));
   AOI22_X1 i_0_314 (.A1(n_0_286), .A2(n_0_211), .B1(n_0_287), .B2(n_0_205), 
      .ZN(n_0_204));
   AOI22_X1 i_0_315 (.A1(n_0_303), .A2(n_0_217), .B1(n_0_302), .B2(n_0_206), 
      .ZN(n_0_205));
   AOI21_X1 i_0_316 (.A(n_0_207), .B1(n_0_306), .B2(n_0_228), .ZN(n_0_206));
   OAI21_X1 i_0_317 (.A(n_0_208), .B1(n_0_306), .B2(n_0_209), .ZN(n_0_207));
   AOI22_X1 i_0_318 (.A1(b[2]), .A2(n_0_305), .B1(b[10]), .B2(n_0_273), .ZN(
      n_0_208));
   NAND2_X1 i_0_319 (.A1(b[18]), .A2(n_0_235), .ZN(n_0_209));
   INV_X1 i_0_320 (.A(n_0_210), .ZN(n_134));
   AOI22_X1 i_0_321 (.A1(n_0_286), .A2(n_0_216), .B1(n_0_287), .B2(n_0_211), 
      .ZN(n_0_210));
   AOI21_X1 i_0_322 (.A(n_0_212), .B1(n_0_303), .B2(n_0_222), .ZN(n_0_211));
   NOR2_X1 i_0_323 (.A1(n_0_303), .A2(n_0_213), .ZN(n_0_212));
   OAI22_X1 i_0_324 (.A1(n_0_306), .A2(n_0_214), .B1(n_0_307), .B2(n_0_234), 
      .ZN(n_0_213));
   AOI222_X1 i_0_325 (.A1(b[19]), .A2(n_0_235), .B1(b[3]), .B2(n_0_308), 
      .C1(b[11]), .C2(n_0_274), .ZN(n_0_214));
   INV_X1 i_0_326 (.A(n_0_215), .ZN(n_135));
   AOI22_X1 i_0_327 (.A1(n_0_286), .A2(n_0_221), .B1(n_0_287), .B2(n_0_216), 
      .ZN(n_0_215));
   AOI22_X1 i_0_328 (.A1(n_0_302), .A2(n_0_217), .B1(n_0_303), .B2(n_0_227), 
      .ZN(n_0_216));
   AOI222_X1 i_0_329 (.A1(b[8]), .A2(n_0_291), .B1(b[16]), .B2(n_0_256), 
      .C1(n_0_307), .C2(n_0_218), .ZN(n_0_217));
   INV_X1 i_0_330 (.A(n_0_219), .ZN(n_0_218));
   AOI222_X1 i_0_331 (.A1(b[20]), .A2(n_0_235), .B1(b[4]), .B2(n_0_308), 
      .C1(b[12]), .C2(n_0_274), .ZN(n_0_219));
   INV_X1 i_0_332 (.A(n_0_220), .ZN(n_136));
   AOI22_X1 i_0_333 (.A1(n_0_286), .A2(n_0_226), .B1(n_0_287), .B2(n_0_221), 
      .ZN(n_0_220));
   AOI22_X1 i_0_334 (.A1(n_0_303), .A2(n_0_232), .B1(n_0_302), .B2(n_0_222), 
      .ZN(n_0_221));
   AOI222_X1 i_0_335 (.A1(b[17]), .A2(n_0_256), .B1(b[9]), .B2(n_0_291), 
      .C1(n_0_307), .C2(n_0_223), .ZN(n_0_222));
   INV_X1 i_0_336 (.A(n_0_224), .ZN(n_0_223));
   AOI222_X1 i_0_337 (.A1(b[13]), .A2(n_0_274), .B1(b[21]), .B2(n_0_235), 
      .C1(b[5]), .C2(n_0_308), .ZN(n_0_224));
   INV_X1 i_0_338 (.A(n_0_225), .ZN(n_137));
   AOI22_X1 i_0_339 (.A1(n_0_286), .A2(n_0_231), .B1(n_0_287), .B2(n_0_226), 
      .ZN(n_0_225));
   AOI22_X1 i_0_340 (.A1(n_0_302), .A2(n_0_227), .B1(n_0_303), .B2(n_0_238), 
      .ZN(n_0_226));
   AOI222_X1 i_0_341 (.A1(b[18]), .A2(n_0_256), .B1(b[10]), .B2(n_0_291), 
      .C1(n_0_307), .C2(n_0_228), .ZN(n_0_227));
   INV_X1 i_0_342 (.A(n_0_229), .ZN(n_0_228));
   AOI222_X1 i_0_343 (.A1(b[6]), .A2(n_0_308), .B1(b[14]), .B2(n_0_274), 
      .C1(b[22]), .C2(n_0_235), .ZN(n_0_229));
   INV_X1 i_0_344 (.A(n_0_230), .ZN(n_138));
   AOI22_X1 i_0_345 (.A1(n_0_286), .A2(n_0_237), .B1(n_0_287), .B2(n_0_231), 
      .ZN(n_0_230));
   AOI22_X1 i_0_346 (.A1(n_0_302), .A2(n_0_232), .B1(n_0_303), .B2(n_0_243), 
      .ZN(n_0_231));
   AOI222_X1 i_0_347 (.A1(b[19]), .A2(n_0_256), .B1(b[11]), .B2(n_0_291), 
      .C1(n_0_307), .C2(n_0_233), .ZN(n_0_232));
   INV_X1 i_0_348 (.A(n_0_234), .ZN(n_0_233));
   AOI222_X1 i_0_349 (.A1(n_155), .A2(n_0_235), .B1(b[7]), .B2(n_0_308), 
      .C1(b[15]), .C2(n_0_274), .ZN(n_0_234));
   AND2_X1 i_0_350 (.A1(n_0_310), .A2(n_0_309), .ZN(n_0_235));
   INV_X1 i_0_351 (.A(n_0_236), .ZN(n_139));
   AOI22_X1 i_0_352 (.A1(n_0_286), .A2(n_0_242), .B1(n_0_287), .B2(n_0_237), 
      .ZN(n_0_236));
   AOI22_X1 i_0_353 (.A1(n_0_302), .A2(n_0_238), .B1(n_0_303), .B2(n_0_248), 
      .ZN(n_0_237));
   AOI221_X1 i_0_354 (.A(n_0_239), .B1(b[20]), .B2(n_0_256), .C1(b[16]), 
      .C2(n_0_273), .ZN(n_0_238));
   INV_X1 i_0_355 (.A(n_0_240), .ZN(n_0_239));
   AOI22_X1 i_0_356 (.A1(b[12]), .A2(n_0_291), .B1(b[8]), .B2(n_0_305), .ZN(
      n_0_240));
   INV_X1 i_0_357 (.A(n_0_241), .ZN(n_140));
   AOI22_X1 i_0_358 (.A1(n_0_286), .A2(n_0_247), .B1(n_0_287), .B2(n_0_242), 
      .ZN(n_0_241));
   AOI22_X1 i_0_359 (.A1(n_0_303), .A2(n_0_253), .B1(n_0_302), .B2(n_0_243), 
      .ZN(n_0_242));
   AOI221_X1 i_0_360 (.A(n_0_244), .B1(b[21]), .B2(n_0_256), .C1(b[17]), 
      .C2(n_0_273), .ZN(n_0_243));
   INV_X1 i_0_361 (.A(n_0_245), .ZN(n_0_244));
   AOI22_X1 i_0_362 (.A1(b[9]), .A2(n_0_305), .B1(b[13]), .B2(n_0_291), .ZN(
      n_0_245));
   INV_X1 i_0_363 (.A(n_0_246), .ZN(n_141));
   AOI22_X1 i_0_364 (.A1(n_0_286), .A2(n_0_252), .B1(n_0_287), .B2(n_0_247), 
      .ZN(n_0_246));
   AOI22_X1 i_0_365 (.A1(n_0_302), .A2(n_0_248), .B1(n_0_303), .B2(n_0_259), 
      .ZN(n_0_247));
   AOI221_X1 i_0_366 (.A(n_0_249), .B1(b[18]), .B2(n_0_273), .C1(b[22]), 
      .C2(n_0_256), .ZN(n_0_248));
   INV_X1 i_0_367 (.A(n_0_250), .ZN(n_0_249));
   AOI22_X1 i_0_368 (.A1(b[14]), .A2(n_0_291), .B1(b[10]), .B2(n_0_305), 
      .ZN(n_0_250));
   INV_X1 i_0_369 (.A(n_0_251), .ZN(n_142));
   AOI22_X1 i_0_370 (.A1(n_0_287), .A2(n_0_252), .B1(n_0_286), .B2(n_0_258), 
      .ZN(n_0_251));
   AOI22_X1 i_0_371 (.A1(n_0_302), .A2(n_0_253), .B1(n_0_303), .B2(n_0_262), 
      .ZN(n_0_252));
   AOI221_X1 i_0_372 (.A(n_0_254), .B1(n_155), .B2(n_0_256), .C1(b[19]), 
      .C2(n_0_273), .ZN(n_0_253));
   INV_X1 i_0_373 (.A(n_0_255), .ZN(n_0_254));
   AOI22_X1 i_0_374 (.A1(b[11]), .A2(n_0_305), .B1(b[15]), .B2(n_0_291), 
      .ZN(n_0_255));
   NOR3_X1 i_0_375 (.A1(n_0_310), .A2(n_0_309), .A3(n_0_307), .ZN(n_0_256));
   INV_X1 i_0_376 (.A(n_0_257), .ZN(n_143));
   AOI22_X1 i_0_377 (.A1(n_0_286), .A2(n_0_261), .B1(n_0_287), .B2(n_0_258), 
      .ZN(n_0_257));
   AOI22_X1 i_0_378 (.A1(n_0_302), .A2(n_0_259), .B1(n_0_303), .B2(n_0_267), 
      .ZN(n_0_258));
   AOI222_X1 i_0_379 (.A1(b[20]), .A2(n_0_273), .B1(b[12]), .B2(n_0_305), 
      .C1(b[16]), .C2(n_0_291), .ZN(n_0_259));
   INV_X1 i_0_380 (.A(n_0_260), .ZN(n_144));
   AOI22_X1 i_0_381 (.A1(n_0_286), .A2(n_0_264), .B1(n_0_287), .B2(n_0_261), 
      .ZN(n_0_260));
   AOI22_X1 i_0_382 (.A1(n_0_302), .A2(n_0_262), .B1(n_0_303), .B2(n_0_272), 
      .ZN(n_0_261));
   AOI222_X1 i_0_383 (.A1(b[21]), .A2(n_0_273), .B1(b[13]), .B2(n_0_305), 
      .C1(b[17]), .C2(n_0_291), .ZN(n_0_262));
   INV_X1 i_0_384 (.A(n_0_263), .ZN(n_145));
   AOI22_X1 i_0_385 (.A1(n_0_287), .A2(n_0_264), .B1(n_0_286), .B2(n_0_269), 
      .ZN(n_0_263));
   OAI21_X1 i_0_386 (.A(n_0_265), .B1(n_0_303), .B2(n_0_267), .ZN(n_0_264));
   AOI21_X1 i_0_387 (.A(n_0_266), .B1(b[16]), .B2(n_0_293), .ZN(n_0_265));
   AND3_X1 i_0_388 (.A1(n_0_303), .A2(n_0_291), .A3(b[20]), .ZN(n_0_266));
   AOI222_X1 i_0_389 (.A1(b[22]), .A2(n_0_273), .B1(b[14]), .B2(n_0_305), 
      .C1(b[18]), .C2(n_0_291), .ZN(n_0_267));
   INV_X1 i_0_390 (.A(n_0_268), .ZN(n_146));
   AOI22_X1 i_0_391 (.A1(n_0_287), .A2(n_0_269), .B1(n_0_286), .B2(n_0_276), 
      .ZN(n_0_268));
   OAI21_X1 i_0_392 (.A(n_0_270), .B1(n_0_303), .B2(n_0_272), .ZN(n_0_269));
   AOI21_X1 i_0_393 (.A(n_0_271), .B1(b[17]), .B2(n_0_293), .ZN(n_0_270));
   AND3_X1 i_0_394 (.A1(n_0_303), .A2(n_0_291), .A3(b[21]), .ZN(n_0_271));
   AOI222_X1 i_0_395 (.A1(n_155), .A2(n_0_273), .B1(b[15]), .B2(n_0_305), 
      .C1(b[19]), .C2(n_0_291), .ZN(n_0_272));
   NOR3_X1 i_0_396 (.A1(n_0_310), .A2(n_0_309), .A3(n_0_306), .ZN(n_0_273));
   NOR2_X1 i_0_397 (.A1(n_0_310), .A2(n_0_309), .ZN(n_0_274));
   INV_X1 i_0_398 (.A(n_0_275), .ZN(n_147));
   AOI22_X1 i_0_399 (.A1(n_0_286), .A2(n_0_279), .B1(n_0_287), .B2(n_0_276), 
      .ZN(n_0_275));
   OAI21_X1 i_0_400 (.A(n_0_277), .B1(n_0_295), .B2(n_0_292), .ZN(n_0_276));
   AOI22_X1 i_0_401 (.A1(b[16]), .A2(n_0_294), .B1(b[18]), .B2(n_0_293), 
      .ZN(n_0_277));
   INV_X1 i_0_402 (.A(n_0_278), .ZN(n_148));
   AOI22_X1 i_0_403 (.A1(n_0_286), .A2(n_0_282), .B1(n_0_287), .B2(n_0_279), 
      .ZN(n_0_278));
   OAI21_X1 i_0_404 (.A(n_0_280), .B1(n_0_297), .B2(n_0_292), .ZN(n_0_279));
   AOI22_X1 i_0_405 (.A1(b[17]), .A2(n_0_294), .B1(b[19]), .B2(n_0_293), 
      .ZN(n_0_280));
   INV_X1 i_0_406 (.A(n_0_281), .ZN(n_149));
   AOI22_X1 i_0_407 (.A1(n_0_288), .A2(n_0_286), .B1(n_0_287), .B2(n_0_282), 
      .ZN(n_0_281));
   OAI21_X1 i_0_408 (.A(n_0_283), .B1(n_0_299), .B2(n_0_292), .ZN(n_0_282));
   AOI22_X1 i_0_409 (.A1(b[18]), .A2(n_0_294), .B1(b[20]), .B2(n_0_293), 
      .ZN(n_0_283));
   INV_X1 i_0_410 (.A(n_0_284), .ZN(n_150));
   AOI21_X1 i_0_411 (.A(n_0_285), .B1(n_0_288), .B2(n_0_287), .ZN(n_0_284));
   NOR3_X1 i_0_412 (.A1(n_0_304), .A2(n_0_295), .A3(n_0_460), .ZN(n_0_285));
   AND2_X1 i_0_413 (.A1(n_0_461), .A2(n_0_312), .ZN(n_0_286));
   AND2_X1 i_0_414 (.A1(n_0_460), .A2(n_0_312), .ZN(n_0_287));
   OAI21_X1 i_0_415 (.A(n_0_289), .B1(n_0_320), .B2(n_0_290), .ZN(n_0_288));
   AOI22_X1 i_0_416 (.A1(b[19]), .A2(n_0_294), .B1(b[21]), .B2(n_0_293), 
      .ZN(n_0_289));
   NAND2_X1 i_0_417 (.A1(n_0_302), .A2(n_0_291), .ZN(n_0_290));
   INV_X1 i_0_418 (.A(n_0_292), .ZN(n_0_291));
   NAND2_X1 i_0_419 (.A1(n_0_308), .A2(n_0_306), .ZN(n_0_292));
   AND2_X1 i_0_420 (.A1(n_0_305), .A2(n_0_303), .ZN(n_0_293));
   AND2_X1 i_0_421 (.A1(n_0_305), .A2(n_0_302), .ZN(n_0_294));
   AOI221_X1 i_0_422 (.A(n_0_304), .B1(n_0_461), .B2(n_0_297), .C1(n_0_460), 
      .C2(n_0_295), .ZN(n_151));
   AOI22_X1 i_0_423 (.A1(b[22]), .A2(n_0_303), .B1(b[20]), .B2(n_0_302), 
      .ZN(n_0_295));
   AOI21_X1 i_0_424 (.A(n_0_304), .B1(n_0_298), .B2(n_0_296), .ZN(n_152));
   OR2_X1 i_0_425 (.A1(n_0_461), .A2(n_0_297), .ZN(n_0_296));
   OAI22_X1 i_0_426 (.A1(b[21]), .A2(n_0_303), .B1(n_155), .B2(n_0_302), 
      .ZN(n_0_297));
   OR2_X1 i_0_427 (.A1(n_0_460), .A2(n_0_299), .ZN(n_0_298));
   NAND2_X1 i_0_428 (.A1(b[22]), .A2(n_0_302), .ZN(n_0_299));
   INV_X1 i_0_429 (.A(n_153), .ZN(n_0_300));
   AOI211_X1 i_0_430 (.A(n_0_301), .B(n_0_304), .C1(n_0_471), .C2(n_0_320), 
      .ZN(n_153));
   OAI21_X1 i_0_431 (.A(n_0_302), .B1(b[22]), .B2(n_0_461), .ZN(n_0_301));
   INV_X1 i_0_432 (.A(n_0_303), .ZN(n_0_302));
   AOI22_X1 i_0_433 (.A1(n_0_467), .A2(n_0_462), .B1(n_0_466), .B2(n_0_463), 
      .ZN(n_0_303));
   NAND2_X1 i_0_434 (.A1(n_0_312), .A2(n_0_305), .ZN(n_0_304));
   NOR3_X1 i_0_435 (.A1(n_0_311), .A2(n_0_309), .A3(n_0_306), .ZN(n_0_305));
   INV_X1 i_0_436 (.A(n_0_307), .ZN(n_0_306));
   XNOR2_X1 i_0_437 (.A(n_0_455), .B(n_0_319), .ZN(n_0_307));
   NOR2_X1 i_0_438 (.A1(n_0_311), .A2(n_0_309), .ZN(n_0_308));
   XNOR2_X1 i_0_439 (.A(n_0_428), .B(n_0_316), .ZN(n_0_309));
   INV_X1 i_0_440 (.A(n_0_311), .ZN(n_0_310));
   OAI21_X1 i_0_441 (.A(n_0_317), .B1(n_0_457), .B2(n_0_318), .ZN(n_0_311));
   AOI21_X1 i_0_442 (.A(n_0_313), .B1(n_0_437), .B2(n_0_315), .ZN(n_0_312));
   AOI211_X1 i_0_443 (.A(n_0_315), .B(n_0_314), .C1(n_0_441), .C2(n_0_439), 
      .ZN(n_0_313));
   AOI211_X1 i_0_444 (.A(n_0_448), .B(n_0_442), .C1(n_0_446), .C2(n_0_443), 
      .ZN(n_0_314));
   OAI21_X1 i_0_445 (.A(n_0_459), .B1(n_0_458), .B2(n_0_316), .ZN(n_0_315));
   OAI21_X1 i_0_446 (.A(n_0_317), .B1(n_0_492), .B2(a[26]), .ZN(n_0_316));
   NAND2_X1 i_0_447 (.A1(n_0_457), .A2(n_0_318), .ZN(n_0_317));
   OAI22_X1 i_0_448 (.A1(n_0_491), .A2(a[25]), .B1(n_0_456), .B2(n_0_319), 
      .ZN(n_0_318));
   AOI21_X1 i_0_449 (.A(n_0_469), .B1(n_0_468), .B2(n_0_462), .ZN(n_0_319));
   NOR2_X1 i_0_450 (.A1(n_0_421), .A2(n_0_320), .ZN(n_154));
   INV_X1 i_0_451 (.A(n_0_320), .ZN(n_155));
   NOR2_X1 i_0_452 (.A1(b[23]), .A2(n_0_475), .ZN(n_0_320));
   OAI22_X1 i_0_453 (.A1(n_0_418), .A2(n_0_325), .B1(n_0_434), .B2(n_0_321), 
      .ZN(n_156));
   AOI22_X1 i_0_454 (.A1(n_0_465), .A2(n_0_322), .B1(n_0_464), .B2(n_0_332), 
      .ZN(n_0_321));
   OAI211_X1 i_0_455 (.A(n_0_324), .B(n_0_323), .C1(n_0_431), .C2(n_0_344), 
      .ZN(n_0_322));
   AOI22_X1 i_0_456 (.A1(a[0]), .A2(n_0_423), .B1(a[8]), .B2(n_0_391), .ZN(
      n_0_323));
   NAND2_X1 i_0_457 (.A1(a[16]), .A2(n_0_339), .ZN(n_0_324));
   OAI21_X1 i_0_458 (.A(n_0_328), .B1(n_0_434), .B2(n_0_325), .ZN(n_157));
   AOI22_X1 i_0_459 (.A1(n_0_465), .A2(n_0_326), .B1(n_0_464), .B2(n_0_337), 
      .ZN(n_0_325));
   AOI22_X1 i_0_460 (.A1(n_0_432), .A2(n_0_349), .B1(n_0_431), .B2(n_0_327), 
      .ZN(n_0_326));
   AOI222_X1 i_0_461 (.A1(a[9]), .A2(n_0_399), .B1(a[1]), .B2(n_0_425), .C1(
      a[17]), .C2(n_0_361), .ZN(n_0_327));
   NAND2_X1 i_0_462 (.A1(n_0_417), .A2(n_0_330), .ZN(n_0_328));
   INV_X1 i_0_463 (.A(n_0_329), .ZN(n_158));
   AOI22_X1 i_0_464 (.A1(n_0_417), .A2(n_0_335), .B1(n_0_433), .B2(n_0_330), 
      .ZN(n_0_329));
   AOI21_X1 i_0_465 (.A(n_0_331), .B1(n_0_464), .B2(n_0_342), .ZN(n_0_330));
   NOR2_X1 i_0_466 (.A1(n_0_464), .A2(n_0_332), .ZN(n_0_331));
   OAI21_X1 i_0_467 (.A(n_0_333), .B1(n_0_431), .B2(n_0_355), .ZN(n_0_332));
   AOI222_X1 i_0_468 (.A1(a[18]), .A2(n_0_339), .B1(a[10]), .B2(n_0_391), 
      .C1(a[2]), .C2(n_0_423), .ZN(n_0_333));
   INV_X1 i_0_469 (.A(n_0_334), .ZN(n_159));
   AOI22_X1 i_0_470 (.A1(n_0_433), .A2(n_0_335), .B1(n_0_417), .B2(n_0_341), 
      .ZN(n_0_334));
   AOI21_X1 i_0_471 (.A(n_0_336), .B1(n_0_464), .B2(n_0_347), .ZN(n_0_335));
   NOR2_X1 i_0_472 (.A1(n_0_464), .A2(n_0_337), .ZN(n_0_336));
   OAI21_X1 i_0_473 (.A(n_0_338), .B1(n_0_431), .B2(n_0_360), .ZN(n_0_337));
   AOI222_X1 i_0_474 (.A1(a[3]), .A2(n_0_423), .B1(a[19]), .B2(n_0_339), 
      .C1(a[11]), .C2(n_0_391), .ZN(n_0_338));
   NOR3_X1 i_0_475 (.A1(n_0_429), .A2(n_0_427), .A3(n_0_432), .ZN(n_0_339));
   INV_X1 i_0_476 (.A(n_0_340), .ZN(n_160));
   AOI22_X1 i_0_477 (.A1(n_0_417), .A2(n_0_346), .B1(n_0_433), .B2(n_0_341), 
      .ZN(n_0_340));
   AOI22_X1 i_0_478 (.A1(n_0_465), .A2(n_0_342), .B1(n_0_464), .B2(n_0_353), 
      .ZN(n_0_341));
   AOI222_X1 i_0_479 (.A1(a[16]), .A2(n_0_378), .B1(a[8]), .B2(n_0_410), 
      .C1(n_0_431), .C2(n_0_343), .ZN(n_0_342));
   INV_X1 i_0_480 (.A(n_0_344), .ZN(n_0_343));
   AOI222_X1 i_0_481 (.A1(a[20]), .A2(n_0_361), .B1(a[12]), .B2(n_0_399), 
      .C1(a[4]), .C2(n_0_425), .ZN(n_0_344));
   INV_X1 i_0_482 (.A(n_0_345), .ZN(n_161));
   AOI22_X1 i_0_483 (.A1(n_0_417), .A2(n_0_351), .B1(n_0_433), .B2(n_0_346), 
      .ZN(n_0_345));
   AOI22_X1 i_0_484 (.A1(n_0_465), .A2(n_0_347), .B1(n_0_464), .B2(n_0_358), 
      .ZN(n_0_346));
   AOI222_X1 i_0_485 (.A1(a[17]), .A2(n_0_378), .B1(a[9]), .B2(n_0_410), 
      .C1(n_0_431), .C2(n_0_348), .ZN(n_0_347));
   INV_X1 i_0_486 (.A(n_0_349), .ZN(n_0_348));
   AOI222_X1 i_0_487 (.A1(a[21]), .A2(n_0_361), .B1(a[13]), .B2(n_0_399), 
      .C1(a[5]), .C2(n_0_425), .ZN(n_0_349));
   INV_X1 i_0_488 (.A(n_0_350), .ZN(n_162));
   AOI22_X1 i_0_489 (.A1(n_0_433), .A2(n_0_351), .B1(n_0_417), .B2(n_0_357), 
      .ZN(n_0_350));
   OAI21_X1 i_0_490 (.A(n_0_352), .B1(n_0_464), .B2(n_0_353), .ZN(n_0_351));
   NAND2_X1 i_0_491 (.A1(n_0_464), .A2(n_0_365), .ZN(n_0_352));
   AOI222_X1 i_0_492 (.A1(a[18]), .A2(n_0_378), .B1(a[10]), .B2(n_0_410), 
      .C1(n_0_431), .C2(n_0_354), .ZN(n_0_353));
   INV_X1 i_0_493 (.A(n_0_355), .ZN(n_0_354));
   AOI222_X1 i_0_494 (.A1(a[22]), .A2(n_0_361), .B1(a[14]), .B2(n_0_399), 
      .C1(a[6]), .C2(n_0_425), .ZN(n_0_355));
   INV_X1 i_0_495 (.A(n_0_356), .ZN(n_163));
   AOI22_X1 i_0_496 (.A1(n_0_417), .A2(n_0_363), .B1(n_0_433), .B2(n_0_357), 
      .ZN(n_0_356));
   AOI22_X1 i_0_497 (.A1(n_0_465), .A2(n_0_358), .B1(n_0_464), .B2(n_0_370), 
      .ZN(n_0_357));
   AOI222_X1 i_0_498 (.A1(a[19]), .A2(n_0_378), .B1(a[11]), .B2(n_0_410), 
      .C1(n_0_431), .C2(n_0_359), .ZN(n_0_358));
   INV_X1 i_0_499 (.A(n_0_360), .ZN(n_0_359));
   AOI222_X1 i_0_500 (.A1(n_180), .A2(n_0_361), .B1(a[15]), .B2(n_0_399), 
      .C1(a[7]), .C2(n_0_425), .ZN(n_0_360));
   NOR2_X1 i_0_501 (.A1(n_0_429), .A2(n_0_427), .ZN(n_0_361));
   INV_X1 i_0_502 (.A(n_0_362), .ZN(n_164));
   AOI22_X1 i_0_503 (.A1(n_0_417), .A2(n_0_369), .B1(n_0_433), .B2(n_0_363), 
      .ZN(n_0_362));
   AOI21_X1 i_0_504 (.A(n_0_364), .B1(n_0_464), .B2(n_0_375), .ZN(n_0_363));
   NOR2_X1 i_0_505 (.A1(n_0_464), .A2(n_0_365), .ZN(n_0_364));
   NAND2_X1 i_0_506 (.A1(n_0_367), .A2(n_0_366), .ZN(n_0_365));
   AOI22_X1 i_0_507 (.A1(a[8]), .A2(n_0_423), .B1(a[12]), .B2(n_0_410), .ZN(
      n_0_366));
   AOI22_X1 i_0_508 (.A1(a[20]), .A2(n_0_378), .B1(a[16]), .B2(n_0_391), 
      .ZN(n_0_367));
   INV_X1 i_0_509 (.A(n_0_368), .ZN(n_165));
   AOI22_X1 i_0_510 (.A1(n_0_417), .A2(n_0_374), .B1(n_0_433), .B2(n_0_369), 
      .ZN(n_0_368));
   AOI22_X1 i_0_511 (.A1(n_0_465), .A2(n_0_370), .B1(n_0_464), .B2(n_0_381), 
      .ZN(n_0_369));
   AOI221_X1 i_0_512 (.A(n_0_371), .B1(a[21]), .B2(n_0_378), .C1(a[17]), 
      .C2(n_0_391), .ZN(n_0_370));
   INV_X1 i_0_513 (.A(n_0_372), .ZN(n_0_371));
   AOI22_X1 i_0_514 (.A1(a[13]), .A2(n_0_410), .B1(a[9]), .B2(n_0_423), .ZN(
      n_0_372));
   INV_X1 i_0_515 (.A(n_0_373), .ZN(n_166));
   AOI22_X1 i_0_516 (.A1(n_0_417), .A2(n_0_380), .B1(n_0_433), .B2(n_0_374), 
      .ZN(n_0_373));
   AOI22_X1 i_0_517 (.A1(n_0_465), .A2(n_0_375), .B1(n_0_464), .B2(n_0_384), 
      .ZN(n_0_374));
   AOI221_X1 i_0_518 (.A(n_0_376), .B1(a[22]), .B2(n_0_378), .C1(a[18]), 
      .C2(n_0_391), .ZN(n_0_375));
   INV_X1 i_0_519 (.A(n_0_377), .ZN(n_0_376));
   AOI22_X1 i_0_520 (.A1(a[14]), .A2(n_0_410), .B1(a[10]), .B2(n_0_423), 
      .ZN(n_0_377));
   NOR3_X1 i_0_521 (.A1(n_0_430), .A2(n_0_426), .A3(n_0_431), .ZN(n_0_378));
   INV_X1 i_0_522 (.A(n_0_379), .ZN(n_167));
   AOI22_X1 i_0_523 (.A1(n_0_417), .A2(n_0_383), .B1(n_0_433), .B2(n_0_380), 
      .ZN(n_0_379));
   AOI22_X1 i_0_524 (.A1(n_0_465), .A2(n_0_381), .B1(n_0_464), .B2(n_0_387), 
      .ZN(n_0_380));
   AOI222_X1 i_0_525 (.A1(a[19]), .A2(n_0_391), .B1(a[11]), .B2(n_0_423), 
      .C1(n_0_432), .C2(n_0_397), .ZN(n_0_381));
   INV_X1 i_0_526 (.A(n_0_382), .ZN(n_168));
   AOI22_X1 i_0_527 (.A1(n_0_417), .A2(n_0_386), .B1(n_0_433), .B2(n_0_383), 
      .ZN(n_0_382));
   AOI22_X1 i_0_528 (.A1(n_0_465), .A2(n_0_384), .B1(n_0_464), .B2(n_0_390), 
      .ZN(n_0_383));
   AOI222_X1 i_0_529 (.A1(a[20]), .A2(n_0_391), .B1(a[12]), .B2(n_0_423), 
      .C1(a[16]), .C2(n_0_410), .ZN(n_0_384));
   INV_X1 i_0_530 (.A(n_0_385), .ZN(n_169));
   AOI22_X1 i_0_531 (.A1(n_0_417), .A2(n_0_389), .B1(n_0_433), .B2(n_0_386), 
      .ZN(n_0_385));
   AOI22_X1 i_0_532 (.A1(n_0_465), .A2(n_0_387), .B1(n_0_464), .B2(n_0_396), 
      .ZN(n_0_386));
   AOI222_X1 i_0_533 (.A1(a[21]), .A2(n_0_391), .B1(a[13]), .B2(n_0_423), 
      .C1(a[17]), .C2(n_0_410), .ZN(n_0_387));
   INV_X1 i_0_534 (.A(n_0_388), .ZN(n_170));
   AOI22_X1 i_0_535 (.A1(n_0_417), .A2(n_0_393), .B1(n_0_433), .B2(n_0_389), 
      .ZN(n_0_388));
   OAI22_X1 i_0_536 (.A1(n_0_465), .A2(n_0_402), .B1(n_0_464), .B2(n_0_390), 
      .ZN(n_0_389));
   AOI222_X1 i_0_537 (.A1(a[22]), .A2(n_0_391), .B1(a[18]), .B2(n_0_410), 
      .C1(a[14]), .C2(n_0_423), .ZN(n_0_390));
   NOR3_X1 i_0_538 (.A1(n_0_430), .A2(n_0_426), .A3(n_0_432), .ZN(n_0_391));
   INV_X1 i_0_539 (.A(n_0_392), .ZN(n_171));
   AOI22_X1 i_0_540 (.A1(n_0_433), .A2(n_0_393), .B1(n_0_417), .B2(n_0_401), 
      .ZN(n_0_392));
   OAI21_X1 i_0_541 (.A(n_0_394), .B1(n_0_464), .B2(n_0_396), .ZN(n_0_393));
   AOI21_X1 i_0_542 (.A(n_0_395), .B1(a[17]), .B2(n_0_411), .ZN(n_0_394));
   AND3_X1 i_0_543 (.A1(a[21]), .A2(n_0_464), .A3(n_0_410), .ZN(n_0_395));
   AOI22_X1 i_0_544 (.A1(a[19]), .A2(n_0_410), .B1(n_0_431), .B2(n_0_397), 
      .ZN(n_0_396));
   INV_X1 i_0_545 (.A(n_0_398), .ZN(n_0_397));
   AOI22_X1 i_0_546 (.A1(n_180), .A2(n_0_399), .B1(a[15]), .B2(n_0_425), 
      .ZN(n_0_398));
   NOR2_X1 i_0_547 (.A1(n_0_430), .A2(n_0_426), .ZN(n_0_399));
   OAI21_X1 i_0_548 (.A(n_0_400), .B1(n_0_418), .B2(n_0_404), .ZN(n_172));
   NAND2_X1 i_0_549 (.A1(n_0_433), .A2(n_0_401), .ZN(n_0_400));
   AOI22_X1 i_0_550 (.A1(n_0_465), .A2(n_0_402), .B1(n_0_464), .B2(n_0_408), 
      .ZN(n_0_401));
   AOI22_X1 i_0_551 (.A1(a[16]), .A2(n_0_423), .B1(a[20]), .B2(n_0_410), 
      .ZN(n_0_402));
   OAI21_X1 i_0_552 (.A(n_0_403), .B1(n_0_434), .B2(n_0_404), .ZN(n_173));
   NAND2_X1 i_0_553 (.A1(n_0_417), .A2(n_0_406), .ZN(n_0_403));
   AOI222_X1 i_0_554 (.A1(n_0_413), .A2(n_0_410), .B1(a[19]), .B2(n_0_411), 
      .C1(a[17]), .C2(n_0_422), .ZN(n_0_404));
   OAI21_X1 i_0_555 (.A(n_0_405), .B1(n_0_418), .B2(n_0_409), .ZN(n_174));
   NAND2_X1 i_0_556 (.A1(n_0_433), .A2(n_0_406), .ZN(n_0_405));
   OAI21_X1 i_0_557 (.A(n_0_407), .B1(n_0_464), .B2(n_0_408), .ZN(n_0_406));
   NAND2_X1 i_0_558 (.A1(a[20]), .A2(n_0_411), .ZN(n_0_407));
   AOI22_X1 i_0_559 (.A1(a[18]), .A2(n_0_423), .B1(a[22]), .B2(n_0_410), 
      .ZN(n_0_408));
   OAI22_X1 i_0_560 (.A1(n_0_434), .A2(n_0_409), .B1(n_0_416), .B2(n_0_412), 
      .ZN(n_175));
   AOI222_X1 i_0_561 (.A1(a[21]), .A2(n_0_411), .B1(n_0_419), .B2(n_0_410), 
      .C1(a[19]), .C2(n_0_422), .ZN(n_0_409));
   NOR3_X1 i_0_562 (.A1(n_0_429), .A2(n_0_426), .A3(n_0_431), .ZN(n_0_410));
   NOR2_X1 i_0_563 (.A1(n_0_465), .A2(n_0_424), .ZN(n_0_411));
   OAI33_X1 i_0_564 (.A1(n_0_434), .A2(n_0_424), .A3(n_0_412), .B1(n_0_424), 
      .B2(n_0_418), .B3(n_0_414), .ZN(n_176));
   AOI22_X1 i_0_565 (.A1(a[22]), .A2(n_0_464), .B1(a[20]), .B2(n_0_465), 
      .ZN(n_0_412));
   OAI33_X1 i_0_566 (.A1(n_0_434), .A2(n_0_424), .A3(n_0_414), .B1(n_0_481), 
      .B2(n_0_464), .B3(n_0_416), .ZN(n_177));
   INV_X1 i_0_567 (.A(n_0_414), .ZN(n_0_413));
   OAI22_X1 i_0_568 (.A1(a[21]), .A2(n_0_464), .B1(n_180), .B2(n_0_465), 
      .ZN(n_0_414));
   OAI21_X1 i_0_569 (.A(n_0_415), .B1(n_0_481), .B2(n_0_421), .ZN(n_178));
   NAND3_X1 i_0_570 (.A1(n_0_423), .A2(n_0_417), .A3(n_0_419), .ZN(n_0_415));
   NAND2_X1 i_0_571 (.A1(n_0_423), .A2(n_0_417), .ZN(n_0_416));
   INV_X1 i_0_572 (.A(n_0_418), .ZN(n_0_417));
   NAND2_X1 i_0_573 (.A1(n_0_461), .A2(n_0_435), .ZN(n_0_418));
   NOR2_X1 i_0_574 (.A1(n_0_477), .A2(n_0_464), .ZN(n_0_419));
   NOR2_X1 i_0_575 (.A1(n_0_477), .A2(n_0_421), .ZN(n_179));
   INV_X1 i_0_576 (.A(n_0_421), .ZN(n_0_420));
   NAND2_X1 i_0_577 (.A1(n_0_433), .A2(n_0_422), .ZN(n_0_421));
   NOR2_X1 i_0_578 (.A1(n_0_464), .A2(n_0_424), .ZN(n_0_422));
   INV_X1 i_0_579 (.A(n_0_424), .ZN(n_0_423));
   NAND2_X1 i_0_580 (.A1(n_0_431), .A2(n_0_425), .ZN(n_0_424));
   NOR2_X1 i_0_581 (.A1(n_0_429), .A2(n_0_426), .ZN(n_0_425));
   INV_X1 i_0_582 (.A(n_0_427), .ZN(n_0_426));
   XNOR2_X1 i_0_583 (.A(n_0_451), .B(n_0_428), .ZN(n_0_427));
   AOI21_X1 i_0_584 (.A(n_0_458), .B1(n_0_493), .B2(a[27]), .ZN(n_0_428));
   INV_X1 i_0_585 (.A(n_0_430), .ZN(n_0_429));
   XNOR2_X1 i_0_586 (.A(n_0_457), .B(n_0_453), .ZN(n_0_430));
   INV_X1 i_0_587 (.A(n_0_432), .ZN(n_0_431));
   XNOR2_X1 i_0_588 (.A(n_0_455), .B(n_0_454), .ZN(n_0_432));
   INV_X1 i_0_589 (.A(n_0_434), .ZN(n_0_433));
   NAND2_X1 i_0_590 (.A1(n_0_460), .A2(n_0_435), .ZN(n_0_434));
   AOI21_X1 i_0_591 (.A(n_0_436), .B1(n_0_449), .B2(n_0_437), .ZN(n_0_435));
   AOI211_X1 i_0_592 (.A(n_0_438), .B(n_0_449), .C1(n_0_447), .C2(n_0_441), 
      .ZN(n_0_436));
   NAND3_X1 i_0_593 (.A1(n_0_441), .A2(n_0_440), .A3(n_0_448), .ZN(n_0_437));
   AOI221_X1 i_0_594 (.A(n_0_440), .B1(n_0_446), .B2(n_0_444), .C1(n_0_445), 
      .C2(n_0_443), .ZN(n_0_438));
   INV_X1 i_0_595 (.A(n_0_440), .ZN(n_0_439));
   NAND2_X1 i_0_596 (.A1(n_0_494), .A2(a[28]), .ZN(n_0_440));
   AND2_X1 i_0_597 (.A1(n_0_446), .A2(n_0_442), .ZN(n_0_441));
   AND2_X1 i_0_598 (.A1(n_0_445), .A2(n_0_444), .ZN(n_0_442));
   INV_X1 i_0_599 (.A(n_0_444), .ZN(n_0_443));
   AOI22_X1 i_0_600 (.A1(b[30]), .A2(n_0_487), .B1(n_0_496), .B2(a[30]), 
      .ZN(n_0_444));
   NAND2_X1 i_0_601 (.A1(n_0_495), .A2(a[29]), .ZN(n_0_445));
   NAND2_X1 i_0_602 (.A1(b[29]), .A2(n_0_486), .ZN(n_0_446));
   INV_X1 i_0_603 (.A(n_0_448), .ZN(n_0_447));
   NAND2_X1 i_0_604 (.A1(b[28]), .A2(n_0_485), .ZN(n_0_448));
   INV_X1 i_0_605 (.A(n_0_450), .ZN(n_0_449));
   AOI21_X1 i_0_606 (.A(n_0_458), .B1(n_0_459), .B2(n_0_451), .ZN(n_0_450));
   AOI22_X1 i_0_607 (.A1(n_0_492), .A2(a[26]), .B1(n_0_457), .B2(n_0_452), 
      .ZN(n_0_451));
   INV_X1 i_0_608 (.A(n_0_453), .ZN(n_0_452));
   AOI21_X1 i_0_609 (.A(n_0_456), .B1(n_0_455), .B2(n_0_454), .ZN(n_0_453));
   AOI21_X1 i_0_610 (.A(n_0_469), .B1(n_0_470), .B2(n_0_468), .ZN(n_0_454));
   AOI21_X1 i_0_611 (.A(n_0_456), .B1(b[25]), .B2(n_0_483), .ZN(n_0_455));
   NOR2_X1 i_0_612 (.A1(b[25]), .A2(n_0_483), .ZN(n_0_456));
   AOI22_X1 i_0_613 (.A1(n_0_492), .A2(a[26]), .B1(b[26]), .B2(n_0_484), 
      .ZN(n_0_457));
   NOR2_X1 i_0_614 (.A1(n_0_493), .A2(a[27]), .ZN(n_0_458));
   NAND2_X1 i_0_615 (.A1(n_0_493), .A2(a[27]), .ZN(n_0_459));
   INV_X1 i_0_616 (.A(n_0_461), .ZN(n_0_460));
   NAND2_X1 i_0_617 (.A1(n_0_470), .A2(n_0_463), .ZN(n_0_461));
   INV_X1 i_0_618 (.A(n_0_463), .ZN(n_0_462));
   NAND2_X1 i_0_619 (.A1(n_0_474), .A2(n_0_471), .ZN(n_0_463));
   INV_X1 i_0_620 (.A(n_0_465), .ZN(n_0_464));
   XNOR2_X1 i_0_621 (.A(n_0_470), .B(n_0_466), .ZN(n_0_465));
   INV_X1 i_0_622 (.A(n_0_467), .ZN(n_0_466));
   OAI21_X1 i_0_623 (.A(n_0_468), .B1(n_0_490), .B2(a[24]), .ZN(n_0_467));
   NAND2_X1 i_0_624 (.A1(n_0_490), .A2(a[24]), .ZN(n_0_468));
   NOR2_X1 i_0_625 (.A1(n_0_490), .A2(a[24]), .ZN(n_0_469));
   NAND2_X1 i_0_626 (.A1(n_0_473), .A2(n_0_472), .ZN(n_0_470));
   INV_X1 i_0_627 (.A(n_0_472), .ZN(n_0_471));
   NAND2_X1 i_0_628 (.A1(n_0_482), .A2(n_0_478), .ZN(n_0_472));
   INV_X1 i_0_629 (.A(n_0_474), .ZN(n_0_473));
   NAND2_X1 i_0_630 (.A1(n_0_489), .A2(n_0_475), .ZN(n_0_474));
   NAND4_X1 i_0_631 (.A1(n_0_495), .A2(n_0_494), .A3(n_0_491), .A4(n_0_476), 
      .ZN(n_0_475));
   NOR4_X1 i_0_632 (.A1(b[26]), .A2(b[24]), .A3(b[30]), .A4(b[27]), .ZN(n_0_476));
   INV_X1 i_0_633 (.A(n_0_477), .ZN(n_180));
   NOR2_X1 i_0_634 (.A1(a[23]), .A2(n_0_478), .ZN(n_0_477));
   NAND4_X1 i_0_635 (.A1(n_0_486), .A2(n_0_485), .A3(n_0_483), .A4(n_0_479), 
      .ZN(n_0_478));
   NOR4_X1 i_0_636 (.A1(a[26]), .A2(a[24]), .A3(a[30]), .A4(a[27]), .ZN(n_0_479));
   INV_X1 i_0_637 (.A(n_0_5), .ZN(n_0_480));
   INV_X1 i_0_638 (.A(a[22]), .ZN(n_0_481));
   INV_X1 i_0_639 (.A(a[23]), .ZN(n_0_482));
   INV_X1 i_0_640 (.A(a[25]), .ZN(n_0_483));
   INV_X1 i_0_641 (.A(a[26]), .ZN(n_0_484));
   INV_X1 i_0_642 (.A(a[28]), .ZN(n_0_485));
   INV_X1 i_0_643 (.A(a[29]), .ZN(n_0_486));
   INV_X1 i_0_644 (.A(a[30]), .ZN(n_0_487));
   INV_X1 i_0_645 (.A(a[31]), .ZN(n_0_488));
   INV_X1 i_0_646 (.A(b[23]), .ZN(n_0_489));
   INV_X1 i_0_647 (.A(b[24]), .ZN(n_0_490));
   INV_X1 i_0_648 (.A(b[25]), .ZN(n_0_491));
   INV_X1 i_0_649 (.A(b[26]), .ZN(n_0_492));
   INV_X1 i_0_650 (.A(b[27]), .ZN(n_0_493));
   INV_X1 i_0_651 (.A(b[28]), .ZN(n_0_494));
   INV_X1 i_0_652 (.A(b[29]), .ZN(n_0_495));
   INV_X1 i_0_653 (.A(b[30]), .ZN(n_0_496));
   INV_X1 i_0_654 (.A(b[31]), .ZN(n_0_497));
   DLH_X1 \i_m_reg[23]  (.D(n_121), .G(n_120), .Q(i_m[23]));
   DLH_X1 \i_m_reg[22]  (.D(n_119), .G(n_120), .Q(i_m[22]));
   DLH_X1 \i_m_reg[21]  (.D(n_118), .G(n_120), .Q(i_m[21]));
   DLH_X1 \i_m_reg[20]  (.D(n_117), .G(n_120), .Q(i_m[20]));
   DLH_X1 \i_m_reg[19]  (.D(n_116), .G(n_120), .Q(i_m[19]));
   DLH_X1 \i_m_reg[18]  (.D(n_115), .G(n_120), .Q(i_m[18]));
   DLH_X1 \i_m_reg[17]  (.D(n_114), .G(n_120), .Q(i_m[17]));
   DLH_X1 \i_m_reg[16]  (.D(n_113), .G(n_120), .Q(i_m[16]));
   DLH_X1 \i_m_reg[15]  (.D(n_112), .G(n_120), .Q(i_m[15]));
   DLH_X1 \i_m_reg[14]  (.D(n_111), .G(n_120), .Q(i_m[14]));
   DLH_X1 \i_m_reg[13]  (.D(n_110), .G(n_120), .Q(i_m[13]));
   DLH_X1 \i_m_reg[12]  (.D(n_109), .G(n_120), .Q(i_m[12]));
   DLH_X1 \i_m_reg[11]  (.D(n_108), .G(n_120), .Q(i_m[11]));
   DLH_X1 \i_m_reg[10]  (.D(n_107), .G(n_120), .Q(i_m[10]));
   DLH_X1 \i_m_reg[9]  (.D(n_106), .G(n_120), .Q(i_m[9]));
   DLH_X1 \i_m_reg[8]  (.D(n_105), .G(n_120), .Q(i_m[8]));
   DLH_X1 \i_m_reg[7]  (.D(n_104), .G(n_120), .Q(i_m[7]));
   DLH_X1 \i_m_reg[6]  (.D(n_103), .G(n_120), .Q(i_m[6]));
   DLH_X1 \i_m_reg[5]  (.D(n_102), .G(n_120), .Q(i_m[5]));
   DLH_X1 \i_m_reg[4]  (.D(n_101), .G(n_120), .Q(i_m[4]));
   DLH_X1 \i_m_reg[3]  (.D(n_100), .G(n_120), .Q(i_m[3]));
   DLH_X1 \i_m_reg[2]  (.D(n_99), .G(n_120), .Q(i_m[2]));
   DLH_X1 \i_m_reg[1]  (.D(n_98), .G(n_120), .Q(i_m[1]));
   DLH_X1 \i_m_reg[0]  (.D(n_97), .G(n_120), .Q(i_m[0]));
   DLH_X1 \i_e_reg[7]  (.D(n_130), .G(n_120), .Q(i_e[7]));
   DLH_X1 \i_e_reg[6]  (.D(n_129), .G(n_120), .Q(i_e[6]));
   DLH_X1 \i_e_reg[5]  (.D(n_128), .G(n_120), .Q(i_e[5]));
   DLH_X1 \i_e_reg[4]  (.D(n_127), .G(n_120), .Q(i_e[4]));
   DLH_X1 \i_e_reg[3]  (.D(n_126), .G(n_120), .Q(i_e[3]));
   DLH_X1 \i_e_reg[2]  (.D(n_125), .G(n_120), .Q(i_e[2]));
   DLH_X1 \i_e_reg[1]  (.D(n_124), .G(n_120), .Q(i_e[1]));
   DLH_X1 \i_e_reg[0]  (.D(n_123), .G(n_120), .Q(i_e[0]));
   DLH_X1 \CSA_IN2_reg[23]  (.D(n_154), .G(n_122), .Q(CSA_IN2[23]));
   DLH_X1 \CSA_IN2_reg[22]  (.D(n_96), .G(n_122), .Q(CSA_IN2[22]));
   DLH_X1 \CSA_IN2_reg[21]  (.D(n_95), .G(n_122), .Q(CSA_IN2[21]));
   DLH_X1 \CSA_IN2_reg[20]  (.D(n_94), .G(n_122), .Q(CSA_IN2[20]));
   DLH_X1 \CSA_IN2_reg[19]  (.D(n_93), .G(n_122), .Q(CSA_IN2[19]));
   DLH_X1 \CSA_IN2_reg[18]  (.D(n_92), .G(n_122), .Q(CSA_IN2[18]));
   DLH_X1 \CSA_IN2_reg[17]  (.D(n_91), .G(n_122), .Q(CSA_IN2[17]));
   DLH_X1 \CSA_IN2_reg[16]  (.D(n_90), .G(n_122), .Q(CSA_IN2[16]));
   DLH_X1 \CSA_IN2_reg[15]  (.D(n_89), .G(n_122), .Q(CSA_IN2[15]));
   DLH_X1 \CSA_IN2_reg[14]  (.D(n_88), .G(n_122), .Q(CSA_IN2[14]));
   DLH_X1 \CSA_IN2_reg[13]  (.D(n_87), .G(n_122), .Q(CSA_IN2[13]));
   DLH_X1 \CSA_IN2_reg[12]  (.D(n_86), .G(n_122), .Q(CSA_IN2[12]));
   DLH_X1 \CSA_IN2_reg[11]  (.D(n_85), .G(n_122), .Q(CSA_IN2[11]));
   DLH_X1 \CSA_IN2_reg[10]  (.D(n_84), .G(n_122), .Q(CSA_IN2[10]));
   DLH_X1 \CSA_IN2_reg[9]  (.D(n_83), .G(n_122), .Q(CSA_IN2[9]));
   DLH_X1 \CSA_IN2_reg[8]  (.D(n_82), .G(n_122), .Q(CSA_IN2[8]));
   DLH_X1 \CSA_IN2_reg[7]  (.D(n_81), .G(n_122), .Q(CSA_IN2[7]));
   DLH_X1 \CSA_IN2_reg[6]  (.D(n_80), .G(n_122), .Q(CSA_IN2[6]));
   DLH_X1 \CSA_IN2_reg[5]  (.D(n_79), .G(n_122), .Q(CSA_IN2[5]));
   DLH_X1 \CSA_IN2_reg[4]  (.D(n_78), .G(n_122), .Q(CSA_IN2[4]));
   DLH_X1 \CSA_IN2_reg[3]  (.D(n_77), .G(n_122), .Q(CSA_IN2[3]));
   DLH_X1 \CSA_IN2_reg[2]  (.D(n_76), .G(n_122), .Q(CSA_IN2[2]));
   DLH_X1 \CSA_IN2_reg[1]  (.D(n_75), .G(n_122), .Q(CSA_IN2[1]));
   DLH_X1 \CSA_IN2_reg[0]  (.D(n_74), .G(n_122), .Q(CSA_IN2[0]));
   DLH_X1 \CSA_IN1_reg[23]  (.D(n_73), .G(n_122), .Q(CSA_IN1[23]));
   DLH_X1 \CSA_IN1_reg[22]  (.D(n_72), .G(n_122), .Q(CSA_IN1[22]));
   DLH_X1 \CSA_IN1_reg[21]  (.D(n_71), .G(n_122), .Q(CSA_IN1[21]));
   DLH_X1 \CSA_IN1_reg[20]  (.D(n_70), .G(n_122), .Q(CSA_IN1[20]));
   DLH_X1 \CSA_IN1_reg[19]  (.D(n_69), .G(n_122), .Q(CSA_IN1[19]));
   DLH_X1 \CSA_IN1_reg[18]  (.D(n_68), .G(n_122), .Q(CSA_IN1[18]));
   DLH_X1 \CSA_IN1_reg[17]  (.D(n_67), .G(n_122), .Q(CSA_IN1[17]));
   DLH_X1 \CSA_IN1_reg[16]  (.D(n_66), .G(n_122), .Q(CSA_IN1[16]));
   DLH_X1 \CSA_IN1_reg[15]  (.D(n_65), .G(n_122), .Q(CSA_IN1[15]));
   DLH_X1 \CSA_IN1_reg[14]  (.D(n_64), .G(n_122), .Q(CSA_IN1[14]));
   DLH_X1 \CSA_IN1_reg[13]  (.D(n_63), .G(n_122), .Q(CSA_IN1[13]));
   DLH_X1 \CSA_IN1_reg[12]  (.D(n_62), .G(n_122), .Q(CSA_IN1[12]));
   DLH_X1 \CSA_IN1_reg[11]  (.D(n_61), .G(n_122), .Q(CSA_IN1[11]));
   DLH_X1 \CSA_IN1_reg[10]  (.D(n_60), .G(n_122), .Q(CSA_IN1[10]));
   DLH_X1 \CSA_IN1_reg[9]  (.D(n_59), .G(n_122), .Q(CSA_IN1[9]));
   DLH_X1 \CSA_IN1_reg[8]  (.D(n_58), .G(n_122), .Q(CSA_IN1[8]));
   DLH_X1 \CSA_IN1_reg[7]  (.D(n_57), .G(n_122), .Q(CSA_IN1[7]));
   DLH_X1 \CSA_IN1_reg[6]  (.D(n_56), .G(n_122), .Q(CSA_IN1[6]));
   DLH_X1 \CSA_IN1_reg[5]  (.D(n_55), .G(n_122), .Q(CSA_IN1[5]));
   DLH_X1 \CSA_IN1_reg[4]  (.D(n_54), .G(n_122), .Q(CSA_IN1[4]));
   DLH_X1 \CSA_IN1_reg[3]  (.D(n_53), .G(n_122), .Q(CSA_IN1[3]));
   DLH_X1 \CSA_IN1_reg[2]  (.D(n_52), .G(n_122), .Q(CSA_IN1[2]));
   DLH_X1 \CSA_IN1_reg[1]  (.D(n_51), .G(n_122), .Q(CSA_IN1[1]));
   DLH_X1 \CSA_IN1_reg[0]  (.D(n_50), .G(n_122), .Q(CSA_IN1[0]));
endmodule

module fpa(A, B, O);
   input [31:0]A;
   input [31:0]B;
   output [31:0]O;

   wire [31:0]adder_out;
   wire [31:0]adder_b_in;
   wire [31:0]adder_a_in;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;

   adder A1 (.a(adder_a_in), .b(adder_b_in), .out(adder_out));
   DLH_X1 \adder_b_in_reg[31]  (.D(B[31]), .G(n_0_0), .Q(adder_b_in[31]));
   DLH_X1 \adder_b_in_reg[30]  (.D(B[30]), .G(n_0_0), .Q(adder_b_in[30]));
   DLH_X1 \adder_b_in_reg[29]  (.D(B[29]), .G(n_0_0), .Q(adder_b_in[29]));
   DLH_X1 \adder_b_in_reg[28]  (.D(B[28]), .G(n_0_0), .Q(adder_b_in[28]));
   DLH_X1 \adder_b_in_reg[27]  (.D(B[27]), .G(n_0_0), .Q(adder_b_in[27]));
   DLH_X1 \adder_b_in_reg[26]  (.D(B[26]), .G(n_0_0), .Q(adder_b_in[26]));
   DLH_X1 \adder_b_in_reg[25]  (.D(B[25]), .G(n_0_0), .Q(adder_b_in[25]));
   DLH_X1 \adder_b_in_reg[24]  (.D(B[24]), .G(n_0_0), .Q(adder_b_in[24]));
   DLH_X1 \adder_b_in_reg[23]  (.D(B[23]), .G(n_0_0), .Q(adder_b_in[23]));
   DLH_X1 \adder_b_in_reg[22]  (.D(B[22]), .G(n_0_0), .Q(adder_b_in[22]));
   DLH_X1 \adder_b_in_reg[21]  (.D(B[21]), .G(n_0_0), .Q(adder_b_in[21]));
   DLH_X1 \adder_b_in_reg[20]  (.D(B[20]), .G(n_0_0), .Q(adder_b_in[20]));
   DLH_X1 \adder_b_in_reg[19]  (.D(B[19]), .G(n_0_0), .Q(adder_b_in[19]));
   DLH_X1 \adder_b_in_reg[18]  (.D(B[18]), .G(n_0_0), .Q(adder_b_in[18]));
   DLH_X1 \adder_b_in_reg[17]  (.D(B[17]), .G(n_0_0), .Q(adder_b_in[17]));
   DLH_X1 \adder_b_in_reg[16]  (.D(B[16]), .G(n_0_0), .Q(adder_b_in[16]));
   DLH_X1 \adder_b_in_reg[15]  (.D(B[15]), .G(n_0_0), .Q(adder_b_in[15]));
   DLH_X1 \adder_b_in_reg[14]  (.D(B[14]), .G(n_0_0), .Q(adder_b_in[14]));
   DLH_X1 \adder_b_in_reg[13]  (.D(B[13]), .G(n_0_0), .Q(adder_b_in[13]));
   DLH_X1 \adder_b_in_reg[12]  (.D(B[12]), .G(n_0_0), .Q(adder_b_in[12]));
   DLH_X1 \adder_b_in_reg[11]  (.D(B[11]), .G(n_0_0), .Q(adder_b_in[11]));
   DLH_X1 \adder_b_in_reg[10]  (.D(B[10]), .G(n_0_0), .Q(adder_b_in[10]));
   DLH_X1 \adder_b_in_reg[9]  (.D(B[9]), .G(n_0_0), .Q(adder_b_in[9]));
   DLH_X1 \adder_b_in_reg[8]  (.D(B[8]), .G(n_0_0), .Q(adder_b_in[8]));
   DLH_X1 \adder_b_in_reg[7]  (.D(B[7]), .G(n_0_0), .Q(adder_b_in[7]));
   DLH_X1 \adder_b_in_reg[6]  (.D(B[6]), .G(n_0_0), .Q(adder_b_in[6]));
   DLH_X1 \adder_b_in_reg[5]  (.D(B[5]), .G(n_0_0), .Q(adder_b_in[5]));
   DLH_X1 \adder_b_in_reg[4]  (.D(B[4]), .G(n_0_0), .Q(adder_b_in[4]));
   DLH_X1 \adder_b_in_reg[3]  (.D(B[3]), .G(n_0_0), .Q(adder_b_in[3]));
   DLH_X1 \adder_b_in_reg[2]  (.D(B[2]), .G(n_0_0), .Q(adder_b_in[2]));
   DLH_X1 \adder_b_in_reg[1]  (.D(B[1]), .G(n_0_0), .Q(adder_b_in[1]));
   DLH_X1 \adder_b_in_reg[0]  (.D(B[0]), .G(n_0_0), .Q(adder_b_in[0]));
   DLH_X1 \adder_a_in_reg[31]  (.D(A[31]), .G(n_0_0), .Q(adder_a_in[31]));
   DLH_X1 \adder_a_in_reg[30]  (.D(A[30]), .G(n_0_0), .Q(adder_a_in[30]));
   DLH_X1 \adder_a_in_reg[29]  (.D(A[29]), .G(n_0_0), .Q(adder_a_in[29]));
   DLH_X1 \adder_a_in_reg[28]  (.D(A[28]), .G(n_0_0), .Q(adder_a_in[28]));
   DLH_X1 \adder_a_in_reg[27]  (.D(A[27]), .G(n_0_0), .Q(adder_a_in[27]));
   DLH_X1 \adder_a_in_reg[26]  (.D(A[26]), .G(n_0_0), .Q(adder_a_in[26]));
   DLH_X1 \adder_a_in_reg[25]  (.D(A[25]), .G(n_0_0), .Q(adder_a_in[25]));
   DLH_X1 \adder_a_in_reg[24]  (.D(A[24]), .G(n_0_0), .Q(adder_a_in[24]));
   DLH_X1 \adder_a_in_reg[23]  (.D(A[23]), .G(n_0_0), .Q(adder_a_in[23]));
   DLH_X1 \adder_a_in_reg[22]  (.D(A[22]), .G(n_0_0), .Q(adder_a_in[22]));
   DLH_X1 \adder_a_in_reg[21]  (.D(A[21]), .G(n_0_0), .Q(adder_a_in[21]));
   DLH_X1 \adder_a_in_reg[20]  (.D(A[20]), .G(n_0_0), .Q(adder_a_in[20]));
   DLH_X1 \adder_a_in_reg[19]  (.D(A[19]), .G(n_0_0), .Q(adder_a_in[19]));
   DLH_X1 \adder_a_in_reg[18]  (.D(A[18]), .G(n_0_0), .Q(adder_a_in[18]));
   DLH_X1 \adder_a_in_reg[17]  (.D(A[17]), .G(n_0_0), .Q(adder_a_in[17]));
   DLH_X1 \adder_a_in_reg[16]  (.D(A[16]), .G(n_0_0), .Q(adder_a_in[16]));
   DLH_X1 \adder_a_in_reg[15]  (.D(A[15]), .G(n_0_0), .Q(adder_a_in[15]));
   DLH_X1 \adder_a_in_reg[14]  (.D(A[14]), .G(n_0_0), .Q(adder_a_in[14]));
   DLH_X1 \adder_a_in_reg[13]  (.D(A[13]), .G(n_0_0), .Q(adder_a_in[13]));
   DLH_X1 \adder_a_in_reg[12]  (.D(A[12]), .G(n_0_0), .Q(adder_a_in[12]));
   DLH_X1 \adder_a_in_reg[11]  (.D(A[11]), .G(n_0_0), .Q(adder_a_in[11]));
   DLH_X1 \adder_a_in_reg[10]  (.D(A[10]), .G(n_0_0), .Q(adder_a_in[10]));
   DLH_X1 \adder_a_in_reg[9]  (.D(A[9]), .G(n_0_0), .Q(adder_a_in[9]));
   DLH_X1 \adder_a_in_reg[8]  (.D(A[8]), .G(n_0_0), .Q(adder_a_in[8]));
   DLH_X1 \adder_a_in_reg[7]  (.D(A[7]), .G(n_0_0), .Q(adder_a_in[7]));
   DLH_X1 \adder_a_in_reg[6]  (.D(A[6]), .G(n_0_0), .Q(adder_a_in[6]));
   DLH_X1 \adder_a_in_reg[5]  (.D(A[5]), .G(n_0_0), .Q(adder_a_in[5]));
   DLH_X1 \adder_a_in_reg[4]  (.D(A[4]), .G(n_0_0), .Q(adder_a_in[4]));
   DLH_X1 \adder_a_in_reg[3]  (.D(A[3]), .G(n_0_0), .Q(adder_a_in[3]));
   DLH_X1 \adder_a_in_reg[2]  (.D(A[2]), .G(n_0_0), .Q(adder_a_in[2]));
   DLH_X1 \adder_a_in_reg[1]  (.D(A[1]), .G(n_0_0), .Q(adder_a_in[1]));
   DLH_X1 \adder_a_in_reg[0]  (.D(A[0]), .G(n_0_0), .Q(adder_a_in[0]));
   INV_X1 i_0_0_0 (.A(n_0_0_0), .ZN(O[0]));
   AOI222_X1 i_0_0_1 (.A1(A[0]), .A2(n_0_0_28), .B1(B[0]), .B2(n_0_0_25), 
      .C1(adder_out[0]), .C2(n_0_0), .ZN(n_0_0_0));
   INV_X1 i_0_0_2 (.A(n_0_0_1), .ZN(O[1]));
   AOI222_X1 i_0_0_3 (.A1(A[1]), .A2(n_0_0_28), .B1(B[1]), .B2(n_0_0_25), 
      .C1(adder_out[1]), .C2(n_0_0), .ZN(n_0_0_1));
   INV_X1 i_0_0_4 (.A(n_0_0_2), .ZN(O[2]));
   AOI222_X1 i_0_0_5 (.A1(A[2]), .A2(n_0_0_28), .B1(B[2]), .B2(n_0_0_25), 
      .C1(adder_out[2]), .C2(n_0_0), .ZN(n_0_0_2));
   INV_X1 i_0_0_6 (.A(n_0_0_3), .ZN(O[3]));
   AOI222_X1 i_0_0_7 (.A1(A[3]), .A2(n_0_0_28), .B1(B[3]), .B2(n_0_0_25), 
      .C1(adder_out[3]), .C2(n_0_0), .ZN(n_0_0_3));
   INV_X1 i_0_0_8 (.A(n_0_0_4), .ZN(O[4]));
   AOI222_X1 i_0_0_9 (.A1(A[4]), .A2(n_0_0_28), .B1(B[4]), .B2(n_0_0_25), 
      .C1(adder_out[4]), .C2(n_0_0), .ZN(n_0_0_4));
   INV_X1 i_0_0_10 (.A(n_0_0_5), .ZN(O[5]));
   AOI222_X1 i_0_0_11 (.A1(A[5]), .A2(n_0_0_28), .B1(B[5]), .B2(n_0_0_25), 
      .C1(adder_out[5]), .C2(n_0_0), .ZN(n_0_0_5));
   INV_X1 i_0_0_12 (.A(n_0_0_6), .ZN(O[6]));
   AOI222_X1 i_0_0_13 (.A1(A[6]), .A2(n_0_0_28), .B1(B[6]), .B2(n_0_0_25), 
      .C1(adder_out[6]), .C2(n_0_0), .ZN(n_0_0_6));
   INV_X1 i_0_0_14 (.A(n_0_0_7), .ZN(O[7]));
   AOI222_X1 i_0_0_15 (.A1(A[7]), .A2(n_0_0_28), .B1(B[7]), .B2(n_0_0_25), 
      .C1(adder_out[7]), .C2(n_0_0), .ZN(n_0_0_7));
   INV_X1 i_0_0_16 (.A(n_0_0_8), .ZN(O[8]));
   AOI222_X1 i_0_0_17 (.A1(A[8]), .A2(n_0_0_28), .B1(B[8]), .B2(n_0_0_25), 
      .C1(adder_out[8]), .C2(n_0_0), .ZN(n_0_0_8));
   INV_X1 i_0_0_18 (.A(n_0_0_9), .ZN(O[9]));
   AOI222_X1 i_0_0_19 (.A1(A[9]), .A2(n_0_0_28), .B1(B[9]), .B2(n_0_0_25), 
      .C1(adder_out[9]), .C2(n_0_0), .ZN(n_0_0_9));
   INV_X1 i_0_0_20 (.A(n_0_0_10), .ZN(O[10]));
   AOI222_X1 i_0_0_21 (.A1(A[10]), .A2(n_0_0_28), .B1(B[10]), .B2(n_0_0_25), 
      .C1(adder_out[10]), .C2(n_0_0), .ZN(n_0_0_10));
   INV_X1 i_0_0_22 (.A(n_0_0_11), .ZN(O[11]));
   AOI222_X1 i_0_0_23 (.A1(A[11]), .A2(n_0_0_28), .B1(B[11]), .B2(n_0_0_25), 
      .C1(adder_out[11]), .C2(n_0_0), .ZN(n_0_0_11));
   INV_X1 i_0_0_24 (.A(n_0_0_12), .ZN(O[12]));
   AOI222_X1 i_0_0_25 (.A1(A[12]), .A2(n_0_0_28), .B1(B[12]), .B2(n_0_0_25), 
      .C1(adder_out[12]), .C2(n_0_0), .ZN(n_0_0_12));
   INV_X1 i_0_0_26 (.A(n_0_0_13), .ZN(O[13]));
   AOI222_X1 i_0_0_27 (.A1(A[13]), .A2(n_0_0_28), .B1(B[13]), .B2(n_0_0_25), 
      .C1(adder_out[13]), .C2(n_0_0), .ZN(n_0_0_13));
   INV_X1 i_0_0_28 (.A(n_0_0_14), .ZN(O[14]));
   AOI222_X1 i_0_0_29 (.A1(A[14]), .A2(n_0_0_28), .B1(B[14]), .B2(n_0_0_25), 
      .C1(adder_out[14]), .C2(n_0_0), .ZN(n_0_0_14));
   INV_X1 i_0_0_30 (.A(n_0_0_15), .ZN(O[15]));
   AOI222_X1 i_0_0_31 (.A1(A[15]), .A2(n_0_0_28), .B1(B[15]), .B2(n_0_0_25), 
      .C1(adder_out[15]), .C2(n_0_0), .ZN(n_0_0_15));
   INV_X1 i_0_0_32 (.A(n_0_0_16), .ZN(O[16]));
   AOI222_X1 i_0_0_33 (.A1(A[16]), .A2(n_0_0_28), .B1(B[16]), .B2(n_0_0_25), 
      .C1(adder_out[16]), .C2(n_0_0), .ZN(n_0_0_16));
   INV_X1 i_0_0_34 (.A(n_0_0_17), .ZN(O[17]));
   AOI222_X1 i_0_0_35 (.A1(A[17]), .A2(n_0_0_28), .B1(B[17]), .B2(n_0_0_25), 
      .C1(adder_out[17]), .C2(n_0_0), .ZN(n_0_0_17));
   INV_X1 i_0_0_36 (.A(n_0_0_18), .ZN(O[18]));
   AOI222_X1 i_0_0_37 (.A1(A[18]), .A2(n_0_0_28), .B1(B[18]), .B2(n_0_0_25), 
      .C1(adder_out[18]), .C2(n_0_0), .ZN(n_0_0_18));
   INV_X1 i_0_0_38 (.A(n_0_0_19), .ZN(O[19]));
   AOI222_X1 i_0_0_39 (.A1(A[19]), .A2(n_0_0_28), .B1(B[19]), .B2(n_0_0_25), 
      .C1(adder_out[19]), .C2(n_0_0), .ZN(n_0_0_19));
   INV_X1 i_0_0_40 (.A(n_0_0_20), .ZN(O[20]));
   AOI222_X1 i_0_0_41 (.A1(A[20]), .A2(n_0_0_28), .B1(B[20]), .B2(n_0_0_25), 
      .C1(adder_out[20]), .C2(n_0_0), .ZN(n_0_0_20));
   INV_X1 i_0_0_42 (.A(n_0_0_21), .ZN(O[21]));
   AOI222_X1 i_0_0_43 (.A1(A[21]), .A2(n_0_0_28), .B1(B[21]), .B2(n_0_0_25), 
      .C1(adder_out[21]), .C2(n_0_0), .ZN(n_0_0_21));
   INV_X1 i_0_0_44 (.A(n_0_0_22), .ZN(O[22]));
   AOI222_X1 i_0_0_45 (.A1(A[22]), .A2(n_0_0_28), .B1(B[22]), .B2(n_0_0_25), 
      .C1(adder_out[22]), .C2(n_0_0), .ZN(n_0_0_22));
   OR2_X1 i_0_0_46 (.A1(adder_out[23]), .A2(n_0_0_24), .ZN(O[23]));
   OR2_X1 i_0_0_47 (.A1(adder_out[24]), .A2(n_0_0_24), .ZN(O[24]));
   OR2_X1 i_0_0_48 (.A1(adder_out[25]), .A2(n_0_0_24), .ZN(O[25]));
   OR2_X1 i_0_0_49 (.A1(adder_out[26]), .A2(n_0_0_24), .ZN(O[26]));
   OR2_X1 i_0_0_50 (.A1(adder_out[27]), .A2(n_0_0_24), .ZN(O[27]));
   OR2_X1 i_0_0_51 (.A1(adder_out[28]), .A2(n_0_0_24), .ZN(O[28]));
   OR2_X1 i_0_0_52 (.A1(adder_out[29]), .A2(n_0_0_24), .ZN(O[29]));
   OR2_X1 i_0_0_53 (.A1(adder_out[30]), .A2(n_0_0_24), .ZN(O[30]));
   INV_X1 i_0_0_54 (.A(n_0_0_23), .ZN(O[31]));
   AOI222_X1 i_0_0_55 (.A1(A[31]), .A2(n_0_0_28), .B1(B[31]), .B2(n_0_0_25), 
      .C1(adder_out[31]), .C2(n_0_0), .ZN(n_0_0_23));
   INV_X1 i_0_0_56 (.A(n_0_0), .ZN(n_0_0_24));
   NOR2_X1 i_0_0_57 (.A1(n_0_0_28), .A2(n_0_0_25), .ZN(n_0_0));
   NOR3_X1 i_0_0_58 (.A1(n_0_0_27), .A2(n_0_0_26), .A3(n_0_0_28), .ZN(n_0_0_25));
   NAND4_X1 i_0_0_59 (.A1(B[30]), .A2(B[29]), .A3(B[28]), .A4(B[27]), .ZN(
      n_0_0_26));
   NAND4_X1 i_0_0_60 (.A1(B[26]), .A2(B[25]), .A3(B[24]), .A4(B[23]), .ZN(
      n_0_0_27));
   NOR2_X1 i_0_0_61 (.A1(n_0_0_30), .A2(n_0_0_29), .ZN(n_0_0_28));
   NAND4_X1 i_0_0_62 (.A1(A[30]), .A2(A[29]), .A3(A[28]), .A4(A[27]), .ZN(
      n_0_0_29));
   NAND4_X1 i_0_0_63 (.A1(A[26]), .A2(A[25]), .A3(A[24]), .A4(A[23]), .ZN(
      n_0_0_30));
endmodule
